magic
tech scmos
timestamp 1525045875
<< metal1 >>
rect 1436 4703 1457 4716
rect 1744 4690 1769 4714
rect 2044 4707 2057 4721
rect 2343 4706 2365 4727
rect 2645 4704 2661 4717
rect 2937 4699 2969 4726
rect 3235 4698 3269 4721
rect 3535 4699 3567 4722
rect 3839 4698 3868 4726
rect 1023 3974 1029 3981
rect 1023 3968 1066 3974
rect 277 3830 307 3868
rect 1060 3729 1066 3968
rect 1323 3959 1329 3981
rect 1623 3960 1629 3981
rect 1923 3960 1929 3981
rect 2223 3960 2229 3981
rect 2523 3960 2529 3981
rect 2907 3976 2992 3990
rect 2919 3968 2979 3976
rect 2931 3960 2970 3968
rect 3123 3960 3129 3981
rect 3423 3960 3429 3981
rect 3723 3960 3729 3981
rect 1622 3959 3729 3960
rect 1323 3958 3729 3959
rect 1323 3953 3962 3958
rect 1123 3935 2107 3943
rect 2331 3920 2783 3929
rect 1090 3907 2050 3916
rect 2315 3884 2908 3893
rect 1019 3723 1066 3729
rect 281 3530 311 3576
rect 1060 3429 1066 3723
rect 2941 3555 2960 3953
rect 3065 3920 3461 3929
rect 3956 3729 3962 3953
rect 4699 3839 4717 3863
rect 3956 3723 3981 3729
rect 2541 3536 2960 3555
rect 4699 3536 4725 3564
rect 1019 3423 1066 3429
rect 275 3229 305 3274
rect 1060 3129 1066 3423
rect 1069 3516 2034 3525
rect 1069 3366 1078 3516
rect 2541 3471 2560 3536
rect 3956 3423 3981 3429
rect 1019 3123 1066 3129
rect 279 2930 301 2971
rect 1060 2829 1066 3123
rect 1019 2823 1066 2829
rect 1011 2690 1030 2696
rect 1011 2677 1044 2690
rect 281 2632 310 2663
rect 1011 2658 1053 2677
rect 1060 2658 1066 2823
rect 3956 3129 3962 3423
rect 4700 3234 4720 3254
rect 3956 3123 3981 3129
rect 3956 2829 3962 3123
rect 4698 2928 4727 2963
rect 3956 2823 3981 2829
rect 1011 2640 1494 2658
rect 1011 2622 1053 2640
rect 1011 2608 1044 2622
rect 1011 2603 1030 2608
rect 1060 2477 1066 2640
rect 1019 2471 1066 2477
rect 1060 1929 1066 2471
rect 3956 2529 3962 2823
rect 4704 2636 4729 2664
rect 3956 2523 3981 2529
rect 3434 2364 3948 2372
rect 3956 2364 3962 2523
rect 3977 2383 3991 2390
rect 3970 2372 3991 2383
rect 3966 2364 3991 2372
rect 3434 2355 3991 2364
rect 3937 2347 3991 2355
rect 3966 2336 3991 2347
rect 3970 2319 3991 2336
rect 4698 2334 4723 2364
rect 3977 2307 3991 2319
rect 4699 2034 4725 2069
rect 1019 1923 1066 1929
rect 3957 1923 3981 1929
rect 277 1726 310 1767
rect 3957 1629 3964 1923
rect 4703 1733 4726 1769
rect 1019 1623 1049 1629
rect 279 1428 306 1474
rect 1042 1329 1049 1623
rect 3957 1623 3981 1629
rect 1019 1323 1049 1329
rect 280 1130 308 1168
rect 1042 1051 1049 1323
rect 2340 1051 2364 1592
rect 3957 1329 3964 1623
rect 4706 1436 4729 1471
rect 3957 1323 3981 1329
rect 3957 1051 3964 1323
rect 4702 1134 4729 1168
rect 1042 1044 3964 1051
rect 1042 1029 1048 1044
rect 1019 1023 1048 1029
rect 1023 1019 1029 1023
rect 1323 1019 1329 1044
rect 1623 1019 1629 1044
rect 1923 1019 1929 1044
rect 2340 1039 2364 1044
rect 2330 1031 2375 1039
rect 2315 1022 2384 1031
rect 2307 1012 2394 1022
rect 2523 1019 2529 1044
rect 2823 1019 2829 1044
rect 3123 1019 3129 1044
rect 3423 1019 3429 1044
rect 3723 1019 3729 1044
rect 3957 1029 3964 1044
rect 3957 1023 3981 1029
rect 1141 280 1166 307
rect 1428 280 1469 305
rect 2033 303 2066 309
rect 1730 280 1764 303
rect 2031 278 2069 303
rect 2325 280 2352 303
rect 2630 276 2669 307
rect 2936 279 2968 304
rect 3224 278 3271 307
rect 3534 284 3566 307
rect 3836 279 3866 308
<< m2contact >>
rect 1023 3981 1029 3987
rect 1323 3981 1329 3987
rect 1623 3981 1629 3987
rect 1923 3981 1929 3987
rect 2223 3981 2229 3987
rect 2523 3981 2529 3987
rect 3123 3981 3129 3987
rect 3423 3981 3429 3987
rect 3723 3981 3729 3987
rect 1115 3935 1123 3943
rect 2107 3935 2115 3943
rect 2322 3920 2331 3929
rect 2783 3920 2793 3929
rect 1081 3907 1090 3916
rect 2050 3907 2059 3916
rect 2306 3884 2315 3893
rect 2908 3884 2917 3893
rect 1013 3723 1019 3729
rect 3055 3920 3065 3929
rect 3461 3920 3470 3929
rect 3981 3723 3987 3729
rect 1013 3423 1019 3429
rect 2034 3516 2043 3525
rect 1069 3357 1078 3366
rect 3981 3423 3987 3429
rect 1013 3123 1019 3129
rect 1013 2823 1019 2829
rect 3981 3123 3987 3129
rect 3981 2823 3987 2829
rect 1494 2640 1512 2658
rect 1013 2471 1019 2477
rect 3981 2523 3987 2529
rect 3417 2355 3434 2372
rect 1013 1923 1019 1929
rect 3981 1923 3987 1929
rect 1013 1623 1019 1629
rect 3981 1623 3987 1629
rect 1013 1323 1019 1329
rect 3981 1323 3987 1329
rect 1013 1023 1019 1029
rect 1023 1013 1029 1019
rect 1323 1013 1329 1019
rect 1623 1013 1629 1019
rect 1923 1013 1929 1019
rect 2523 1013 2529 1019
rect 2823 1013 2829 1019
rect 3123 1013 3129 1019
rect 3423 1013 3429 1019
rect 3981 1023 3987 1029
rect 3723 1013 3729 1019
<< metal2 >>
rect 1346 3975 1351 3984
rect 1346 3970 1408 3975
rect 1647 3970 1652 3984
rect 1945 3978 1952 3984
rect 2245 3974 2252 3985
rect 1019 3957 1032 3966
rect 1024 3943 1032 3957
rect 1024 3935 1115 3943
rect 1081 3666 1090 3907
rect 1018 3657 1090 3666
rect 1019 3357 1069 3366
rect 1014 3058 1036 3065
rect 1403 2720 1408 3970
rect 1420 3965 1652 3970
rect 1420 2790 1425 3965
rect 2549 3950 2553 3985
rect 1975 3946 2553 3950
rect 1430 3898 1484 3903
rect 1430 3284 1435 3898
rect 1438 3886 1528 3891
rect 1438 3292 1443 3886
rect 1975 3500 1979 3946
rect 3149 3943 3153 3985
rect 2039 3500 2043 3516
rect 2055 3500 2059 3907
rect 2111 3500 2115 3935
rect 2279 3939 3153 3943
rect 2279 3500 2283 3939
rect 3449 3936 3453 3985
rect 3745 3976 3750 3981
rect 2343 3932 3453 3936
rect 2311 3503 2315 3884
rect 2311 3502 2314 3503
rect 2327 3500 2331 3920
rect 2343 3500 2347 3932
rect 2793 3920 3055 3929
rect 3470 3920 3953 3929
rect 2423 3908 3940 3917
rect 2423 3500 2427 3908
rect 2879 3896 3928 3905
rect 2879 3500 2883 3896
rect 2917 3884 3916 3893
rect 3907 3629 3916 3884
rect 3919 3641 3928 3896
rect 3931 3653 3940 3908
rect 3944 3666 3953 3920
rect 3978 3746 3983 3751
rect 3944 3657 3981 3666
rect 3931 3644 3953 3653
rect 3919 3632 3941 3641
rect 3907 3620 3929 3629
rect 3920 3342 3929 3620
rect 3932 3354 3941 3632
rect 3944 3366 3953 3644
rect 3944 3357 3981 3366
rect 3932 3345 3953 3354
rect 3920 3333 3941 3342
rect 1438 3287 1448 3292
rect 1430 3279 1439 3284
rect 1434 2848 1439 3279
rect 1443 2860 1448 3287
rect 3932 3054 3941 3333
rect 3944 3066 3953 3345
rect 3944 3057 3981 3066
rect 3932 3045 3953 3054
rect 1434 2843 1450 2848
rect 1445 2814 1450 2843
rect 3944 2766 3953 3045
rect 3944 2757 3981 2766
rect 3964 1945 3984 1952
rect 1016 1647 1061 1650
rect 1016 1347 1055 1350
rect 1052 1087 1055 1347
rect 1058 1093 1061 1647
rect 3975 1645 3985 1652
rect 2536 1093 2539 1563
rect 1058 1090 2539 1093
rect 2552 1087 2555 1564
rect 1052 1084 2555 1087
rect 2640 1081 2643 1563
rect 1019 1078 2643 1081
rect 1019 1044 1022 1078
rect 2656 1075 2659 1563
rect 1103 1072 2659 1075
rect 1103 1018 1106 1072
rect 2672 1069 2675 1563
rect 1346 1066 2675 1069
rect 1049 1015 1106 1018
rect 1346 1016 1349 1066
rect 2704 1063 2707 1564
rect 1646 1060 2707 1063
rect 1646 1016 1649 1060
rect 2720 1057 2723 1563
rect 1944 1054 2723 1057
rect 1944 1013 1947 1054
rect 2736 1036 2739 1563
rect 2816 1061 2819 1565
rect 3976 1345 3986 1352
rect 2816 1058 2850 1061
rect 2544 1033 2739 1036
rect 2544 1013 2547 1033
rect 2847 1014 2850 1058
rect 3978 1045 3986 1052
rect 3145 1016 3152 1023
rect 3745 1028 3752 1031
rect 3445 1016 3452 1023
rect 3744 1019 3753 1028
<< m3contact >>
rect 1945 3971 1952 3978
rect 1036 3058 1043 3065
rect 2245 3967 2252 3974
rect 1484 3898 1489 3903
rect 1528 3886 1533 3891
rect 3745 3971 3750 3976
rect 3973 3746 3978 3751
rect 1443 2855 1448 2860
rect 1445 2809 1450 2814
rect 1420 2785 1425 2790
rect 1403 2715 1408 2720
rect 3957 1945 3964 1952
rect 3968 1645 3975 1652
rect 3969 1345 3976 1352
rect 3971 1045 3978 1052
rect 3745 1031 3752 1038
rect 3145 1023 3152 1030
rect 3445 1023 3452 1030
<< metal3 >>
rect 1944 3978 1953 3979
rect 1944 3971 1945 3978
rect 1952 3971 1953 3978
rect 3744 3976 3751 3977
rect 1944 3970 1953 3971
rect 1948 3932 1953 3970
rect 2244 3974 2253 3975
rect 2244 3967 2245 3974
rect 2252 3967 2253 3974
rect 3744 3971 3745 3976
rect 3750 3971 3751 3976
rect 3744 3970 3751 3971
rect 2244 3966 2253 3967
rect 1446 3927 1953 3932
rect 1446 3300 1451 3927
rect 2248 3924 2253 3966
rect 1454 3919 2253 3924
rect 1454 3380 1459 3919
rect 3745 3913 3750 3970
rect 2271 3908 3750 3913
rect 1483 3903 1490 3904
rect 2271 3903 2276 3908
rect 1483 3898 1484 3903
rect 1489 3898 2276 3903
rect 1483 3897 1490 3898
rect 2291 3896 3978 3901
rect 1527 3891 1534 3892
rect 2291 3891 2296 3896
rect 1527 3886 1528 3891
rect 1533 3886 2296 3891
rect 1527 3885 1534 3886
rect 3973 3752 3978 3896
rect 3972 3751 3979 3752
rect 3972 3746 3973 3751
rect 3978 3746 3979 3751
rect 3972 3745 3979 3746
rect 1446 3295 1454 3300
rect 1035 3065 1044 3066
rect 1035 3058 1036 3065
rect 1043 3058 1044 3065
rect 1035 3057 1044 3058
rect 1039 2900 1044 3057
rect 1039 2895 1454 2900
rect 1442 2860 1449 2861
rect 1442 2855 1443 2860
rect 1448 2855 1454 2860
rect 1442 2854 1449 2855
rect 1444 2814 1451 2815
rect 1454 2814 1459 2815
rect 1444 2809 1445 2814
rect 1450 2809 1459 2814
rect 1444 2808 1451 2809
rect 1419 2790 1426 2791
rect 1419 2785 1420 2790
rect 1425 2785 1454 2790
rect 1419 2784 1426 2785
rect 1402 2720 1409 2721
rect 1402 2715 1403 2720
rect 1408 2715 1454 2720
rect 1402 2714 1409 2715
rect 3474 2345 3932 2350
rect 3927 2342 3932 2345
rect 3927 2337 3961 2342
rect 3474 2325 3952 2330
rect 3474 2275 3943 2280
rect 3474 2255 3935 2260
rect 3474 2235 3927 2240
rect 3474 2165 3919 2170
rect 3474 2135 3911 2140
rect 3906 1075 3911 2135
rect 3144 1070 3911 1075
rect 3144 1030 3153 1070
rect 3914 1067 3919 2165
rect 3144 1023 3145 1030
rect 3152 1023 3153 1030
rect 3144 1022 3153 1023
rect 3444 1062 3919 1067
rect 3444 1030 3453 1062
rect 3922 1059 3927 2235
rect 3745 1054 3927 1059
rect 3745 1039 3752 1054
rect 3930 1051 3935 2255
rect 3938 1349 3943 2275
rect 3947 1649 3952 2325
rect 3956 1953 3961 2337
rect 3956 1952 3965 1953
rect 3956 1945 3957 1952
rect 3964 1945 3965 1952
rect 3956 1944 3965 1945
rect 3967 1652 3976 1653
rect 3967 1649 3968 1652
rect 3947 1645 3968 1649
rect 3975 1645 3976 1652
rect 3947 1644 3976 1645
rect 3968 1352 3977 1353
rect 3968 1349 3969 1352
rect 3938 1345 3969 1349
rect 3976 1345 3977 1352
rect 3938 1344 3977 1345
rect 3970 1052 3979 1053
rect 3970 1051 3971 1052
rect 3930 1046 3971 1051
rect 3970 1045 3971 1046
rect 3978 1045 3979 1052
rect 3970 1044 3979 1045
rect 3744 1038 3753 1039
rect 3744 1031 3745 1038
rect 3752 1031 3753 1038
rect 3744 1030 3753 1031
rect 3444 1023 3445 1030
rect 3452 1023 3453 1030
rect 3444 1022 3453 1023
rect 3445 1016 3452 1022
use top_module  top_module_0
timestamp 1524952243
transform 1 0 1454 0 1 1563
box 0 0 2020 1940
use PadFrame  PadFrame_0
timestamp 1524078036
transform 1 0 2500 0 1 2500
box -2500 -2500 2500 2500
<< labels >>
rlabel metal1 2050 4714 2050 4714 1 p_out_win
rlabel metal1 2352 4715 2352 4715 1 p_out_lose
rlabel metal1 2652 4710 2652 4710 1 p_out_state[1]
rlabel metal1 2953 4712 2953 4712 1 Vdd
rlabel metal1 3247 4708 3247 4708 1 p_out_state[0]
rlabel metal1 3550 4711 3550 4711 1 p_out_state[2]
rlabel metal1 4711 3553 4711 3553 1 p_in_wai
rlabel metal1 4710 3241 4710 3241 1 p_in_clkb
rlabel metal1 4717 2945 4717 2945 1 p_in_clka
rlabel metal1 4717 2650 4717 2650 1 p_in_reset
rlabel metal1 4710 2344 4710 2344 1 Gnd
rlabel metal1 4717 1749 4717 1749 1 p_out_MuxData[0]
rlabel metal1 4708 2051 4708 2051 1 p_out_MuxData[1]
rlabel metal1 4717 1449 4717 1449 1 p_out_MuxData[2]
rlabel metal1 4715 1152 4715 1152 1 p_out_MuxData[3]
rlabel metal1 3854 295 3854 295 1 p_out_MuxData[8]
rlabel metal1 3554 297 3554 297 1 p_out_MuxData[9]
rlabel metal1 3252 297 3252 297 1 p_out_MuxData[10]
rlabel metal1 2951 290 2951 290 1 p_out_MuxData[11]
rlabel metal1 2651 291 2651 291 1 p_out_MuxData[5]
rlabel metal1 2341 291 2341 291 1 Vdd
rlabel metal1 2052 289 2052 289 1 p_out_MuxData[13]
rlabel metal1 1749 288 1749 288 1 p_out_MuxData[15]
rlabel metal1 1448 291 1448 291 1 p_out_MuxData[14]
rlabel metal1 1156 287 1156 287 1 p_out_MuxData[7]
rlabel metal1 297 1153 297 1153 1 p_out_MuxData[6]
rlabel metal1 291 1453 291 1453 1 p_out_MuxData[4]
rlabel metal1 290 1752 290 1752 1 p_out_MuxData[12]
rlabel metal1 294 2646 294 2646 1 Gnd
rlabel metal1 290 2953 290 2953 1 p_in_DataIn
rlabel metal1 291 3253 291 3253 1 p_in_run
rlabel metal1 301 3554 301 3554 1 p_in_timer5
rlabel metal1 293 3852 293 3852 1 p_in_inp
rlabel metal1 4707 3850 4707 3850 1 p_con_count[1]
rlabel metal1 3851 4712 3851 4712 1 p_con_count[3]
rlabel metal1 1758 4703 1758 4703 1 p_con_count[0]
rlabel metal1 1447 4710 1447 4710 1 p_con_count[2]
<< end >>
