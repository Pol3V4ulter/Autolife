magic
tech scmos
timestamp 1524952243
<< metal1 >>
rect 14 1907 2004 1927
rect 38 1883 1980 1903
rect 14 1867 2004 1873
rect 330 1833 348 1836
rect 796 1833 805 1836
rect 898 1833 908 1836
rect 186 1816 189 1825
rect 834 1816 837 1825
rect 186 1813 196 1816
rect 276 1813 293 1816
rect 306 1813 316 1816
rect 402 1813 420 1816
rect 492 1813 509 1816
rect 564 1813 573 1816
rect 588 1813 604 1816
rect 644 1813 653 1816
rect 700 1813 709 1816
rect 772 1813 781 1816
rect 826 1813 837 1816
rect 1074 1813 1092 1816
rect 1164 1813 1181 1816
rect 1234 1813 1244 1816
rect 1300 1813 1308 1816
rect 1386 1813 1396 1816
rect 1428 1813 1437 1816
rect 1580 1813 1597 1816
rect 1636 1813 1644 1816
rect 1676 1813 1685 1816
rect 1738 1813 1756 1816
rect 1828 1813 1837 1816
rect 284 1803 292 1806
rect 580 1803 589 1806
rect 610 1803 620 1806
rect 636 1803 645 1806
rect 650 1805 653 1813
rect 682 1803 692 1806
rect 706 1805 709 1813
rect 826 1805 829 1813
rect 876 1803 885 1806
rect 1236 1803 1245 1806
rect 1274 1803 1285 1806
rect 1292 1803 1301 1806
rect 1370 1803 1380 1806
rect 1282 1795 1285 1803
rect 1386 1795 1389 1813
rect 1394 1803 1404 1806
rect 1426 1803 1436 1806
rect 1674 1803 1684 1806
rect 1826 1803 1836 1806
rect 38 1767 1980 1773
rect 298 1733 308 1736
rect 604 1733 613 1736
rect 852 1733 861 1736
rect 876 1733 900 1736
rect 906 1733 924 1736
rect 1268 1733 1277 1736
rect 1668 1733 1677 1736
rect 1908 1733 1933 1736
rect 826 1726 829 1733
rect 66 1723 76 1726
rect 180 1723 189 1726
rect 452 1723 485 1726
rect 500 1723 517 1726
rect 554 1723 564 1726
rect 578 1723 588 1726
rect 762 1723 772 1726
rect 820 1723 829 1726
rect 850 1723 860 1726
rect 906 1725 909 1733
rect 1010 1726 1013 1733
rect 940 1723 949 1726
rect 988 1723 997 1726
rect 1004 1723 1013 1726
rect 1074 1723 1092 1726
rect 1180 1723 1197 1726
rect 234 1713 244 1716
rect 850 1715 853 1723
rect 946 1715 949 1723
rect 1274 1716 1277 1733
rect 1340 1723 1349 1726
rect 1516 1723 1533 1726
rect 1674 1716 1677 1733
rect 1740 1723 1749 1726
rect 1772 1723 1788 1726
rect 1274 1713 1284 1716
rect 1314 1713 1324 1716
rect 1450 1713 1460 1716
rect 1490 1713 1500 1716
rect 1596 1713 1605 1716
rect 1674 1713 1684 1716
rect 1714 1713 1724 1716
rect 1738 1713 1756 1716
rect 14 1667 2004 1673
rect 386 1616 389 1625
rect 402 1623 436 1626
rect 1250 1623 1260 1626
rect 1786 1623 1796 1626
rect 66 1613 76 1616
rect 322 1613 333 1616
rect 340 1613 357 1616
rect 364 1613 389 1616
rect 396 1613 413 1616
rect 444 1613 461 1616
rect 674 1613 692 1616
rect 828 1613 837 1616
rect 866 1613 876 1616
rect 322 1607 325 1613
rect 354 1607 357 1613
rect 914 1607 917 1616
rect 980 1613 988 1616
rect 994 1613 1004 1616
rect 1092 1613 1109 1616
rect 1162 1613 1172 1616
rect 1204 1613 1213 1616
rect 1276 1613 1285 1616
rect 1548 1613 1565 1616
rect 1612 1613 1621 1616
rect 1692 1613 1709 1616
rect 1786 1606 1789 1623
rect 1858 1613 1876 1616
rect 404 1603 437 1606
rect 452 1603 460 1606
rect 820 1603 836 1606
rect 866 1603 884 1606
rect 1020 1603 1028 1606
rect 1164 1603 1173 1606
rect 1780 1603 1789 1606
rect 866 1595 869 1603
rect 38 1567 1980 1573
rect 708 1543 717 1546
rect 266 1526 269 1534
rect 290 1533 300 1536
rect 66 1523 76 1526
rect 204 1523 221 1526
rect 260 1523 269 1526
rect 314 1523 317 1534
rect 338 1523 356 1526
rect 370 1523 373 1534
rect 394 1523 397 1534
rect 402 1523 405 1534
rect 530 1523 533 1534
rect 682 1533 692 1536
rect 724 1533 733 1536
rect 1058 1533 1068 1536
rect 1090 1533 1100 1536
rect 1588 1533 1597 1536
rect 1730 1533 1740 1536
rect 1818 1533 1828 1536
rect 540 1523 557 1526
rect 708 1523 716 1526
rect 778 1523 796 1526
rect 874 1523 892 1526
rect 930 1523 940 1526
rect 1092 1523 1101 1526
rect 1586 1523 1596 1526
rect 1724 1523 1732 1526
rect 1770 1523 1780 1526
rect 1820 1523 1829 1526
rect 1836 1523 1845 1526
rect 554 1515 557 1523
rect 14 1467 2004 1473
rect 394 1416 397 1425
rect 826 1416 829 1425
rect 74 1413 84 1416
rect 188 1413 197 1416
rect 252 1413 261 1416
rect 282 1405 285 1416
rect 378 1413 388 1416
rect 394 1413 405 1416
rect 412 1413 421 1416
rect 434 1413 444 1416
rect 522 1413 540 1416
rect 564 1413 573 1416
rect 818 1413 829 1416
rect 338 1403 348 1406
rect 394 1403 404 1406
rect 524 1403 533 1406
rect 780 1403 796 1406
rect 818 1405 821 1413
rect 978 1406 981 1414
rect 972 1403 981 1406
rect 1010 1403 1013 1414
rect 1122 1405 1125 1416
rect 1210 1413 1220 1416
rect 1298 1413 1308 1416
rect 1156 1403 1164 1406
rect 1210 1405 1213 1413
rect 1338 1406 1341 1414
rect 1444 1413 1453 1416
rect 1596 1413 1605 1416
rect 1650 1413 1660 1416
rect 1306 1403 1316 1406
rect 1338 1403 1349 1406
rect 1450 1405 1453 1413
rect 1562 1403 1572 1406
rect 1588 1403 1597 1406
rect 1650 1405 1653 1413
rect 1690 1405 1693 1416
rect 1884 1413 1893 1416
rect 1890 1405 1893 1413
rect 338 1395 341 1403
rect 38 1367 1980 1373
rect 170 1336 173 1345
rect 146 1333 173 1336
rect 194 1326 197 1336
rect 228 1333 236 1336
rect 84 1323 101 1326
rect 122 1323 140 1326
rect 194 1325 205 1326
rect 196 1323 205 1325
rect 282 1323 292 1326
rect 298 1323 301 1334
rect 394 1323 404 1326
rect 442 1323 445 1334
rect 724 1333 740 1336
rect 780 1333 796 1336
rect 452 1323 461 1326
rect 514 1323 524 1326
rect 676 1323 685 1326
rect 826 1323 836 1326
rect 954 1325 957 1336
rect 986 1333 996 1336
rect 1106 1323 1116 1326
rect 1146 1323 1155 1326
rect 1210 1323 1213 1333
rect 1258 1323 1261 1334
rect 1348 1333 1357 1336
rect 1380 1333 1389 1336
rect 1514 1326 1517 1336
rect 1546 1333 1564 1336
rect 1586 1326 1589 1336
rect 1610 1333 1620 1336
rect 1666 1326 1669 1336
rect 1292 1323 1317 1326
rect 1410 1323 1420 1326
rect 1474 1323 1492 1326
rect 1594 1323 1602 1326
rect 1618 1323 1627 1326
rect 1682 1323 1685 1334
rect 1730 1323 1733 1334
rect 1786 1323 1789 1334
rect 1908 1333 1916 1336
rect 1900 1323 1924 1326
rect 98 1315 101 1323
rect 316 1313 325 1316
rect 1172 1313 1180 1316
rect 1876 1313 1884 1316
rect 314 1303 332 1306
rect 1660 1303 1669 1306
rect 14 1267 2004 1273
rect 180 1233 197 1236
rect 1434 1233 1452 1236
rect 186 1223 196 1226
rect 394 1216 397 1225
rect 1410 1223 1436 1226
rect 1482 1216 1485 1225
rect 66 1213 76 1216
rect 114 1213 132 1216
rect 244 1213 252 1216
rect 356 1213 373 1216
rect 394 1213 412 1216
rect 468 1213 484 1216
rect 202 1203 212 1206
rect 236 1203 245 1206
rect 250 1203 260 1206
rect 314 1203 324 1206
rect 370 1205 373 1213
rect 466 1203 476 1206
rect 498 1205 501 1216
rect 516 1213 533 1216
rect 546 1213 556 1216
rect 578 1206 581 1214
rect 612 1213 621 1216
rect 628 1213 637 1216
rect 690 1213 708 1216
rect 524 1203 532 1206
rect 572 1203 581 1206
rect 610 1203 620 1206
rect 842 1205 845 1216
rect 914 1213 924 1216
rect 954 1206 957 1215
rect 906 1203 916 1206
rect 948 1203 957 1206
rect 986 1203 996 1206
rect 1106 1205 1109 1216
rect 1122 1205 1125 1216
rect 1132 1213 1141 1216
rect 1154 1205 1157 1216
rect 1330 1205 1333 1216
rect 1466 1213 1476 1216
rect 1482 1213 1492 1216
rect 1498 1213 1508 1216
rect 1412 1203 1429 1206
rect 1498 1205 1501 1213
rect 1538 1206 1541 1214
rect 1610 1213 1627 1216
rect 1666 1213 1676 1216
rect 1698 1213 1708 1216
rect 1746 1213 1756 1216
rect 1844 1213 1885 1216
rect 1932 1213 1941 1216
rect 1524 1203 1541 1206
rect 1706 1203 1716 1206
rect 1940 1203 1949 1206
rect 38 1167 1980 1173
rect 314 1133 324 1136
rect 396 1133 412 1136
rect 524 1133 533 1136
rect 666 1126 669 1135
rect 754 1126 757 1135
rect 796 1133 812 1136
rect 1314 1133 1324 1136
rect 1450 1126 1453 1135
rect 188 1123 212 1126
rect 410 1123 429 1126
rect 452 1123 461 1126
rect 468 1123 485 1126
rect 516 1123 525 1126
rect 540 1123 549 1126
rect 588 1123 605 1126
rect 660 1123 669 1126
rect 716 1123 725 1126
rect 746 1123 757 1126
rect 810 1123 820 1126
rect 988 1123 997 1126
rect 1036 1123 1053 1126
rect 1092 1123 1101 1126
rect 1178 1123 1188 1126
rect 1444 1123 1453 1126
rect 1498 1126 1501 1135
rect 1506 1133 1516 1136
rect 1538 1133 1547 1136
rect 1596 1133 1605 1136
rect 1634 1133 1644 1136
rect 1748 1133 1757 1136
rect 1844 1133 1853 1136
rect 1498 1123 1508 1126
rect 1538 1125 1541 1133
rect 1546 1123 1564 1126
rect 1636 1123 1645 1126
rect 1732 1123 1749 1126
rect 1754 1125 1757 1133
rect 1828 1123 1845 1126
rect 1906 1123 1916 1126
rect 500 1113 508 1116
rect 746 1115 749 1123
rect 14 1067 2004 1073
rect 194 1016 197 1025
rect 1002 1016 1005 1026
rect 1234 1016 1237 1025
rect 66 1013 76 1016
rect 180 1013 197 1016
rect 260 1013 269 1016
rect 354 1006 357 1014
rect 484 1013 493 1016
rect 540 1013 557 1016
rect 762 1014 772 1016
rect 762 1013 773 1014
rect 186 1003 196 1006
rect 245 1003 252 1006
rect 290 1003 308 1006
rect 348 1003 357 1006
rect 380 1003 389 1006
rect 490 1005 493 1013
rect 770 1003 773 1013
rect 1002 1013 1020 1016
rect 1138 1013 1156 1016
rect 1170 1013 1188 1016
rect 1210 1013 1220 1016
rect 1234 1013 1252 1016
rect 1292 1013 1325 1016
rect 1420 1013 1429 1016
rect 1442 1013 1453 1016
rect 804 1003 820 1006
rect 876 1003 885 1006
rect 914 1003 924 1006
rect 1002 1005 1005 1013
rect 1258 1003 1268 1006
rect 1322 1005 1325 1013
rect 1450 1005 1453 1013
rect 1498 1005 1501 1016
rect 1506 1013 1516 1016
rect 1570 1013 1580 1016
rect 1634 1013 1652 1016
rect 1682 1013 1693 1016
rect 1570 1005 1573 1013
rect 1578 1003 1588 1006
rect 1604 1003 1613 1006
rect 1690 1005 1693 1013
rect 1746 1006 1749 1014
rect 1812 1013 1845 1016
rect 1876 1013 1900 1016
rect 1740 1003 1749 1006
rect 1772 1003 1788 1006
rect 1892 1003 1901 1006
rect 1924 1003 1949 1006
rect 292 993 301 996
rect 788 993 796 996
rect 38 967 1980 973
rect 202 926 205 934
rect 194 923 205 926
rect 282 923 285 934
rect 308 933 324 936
rect 330 933 340 936
rect 386 933 396 936
rect 506 926 509 934
rect 882 926 885 934
rect 956 933 965 936
rect 972 933 988 936
rect 332 923 348 926
rect 500 923 509 926
rect 556 923 573 926
rect 748 923 757 926
rect 804 923 821 926
rect 874 923 885 926
rect 1034 923 1037 934
rect 1058 923 1061 934
rect 1106 926 1109 934
rect 1106 923 1116 926
rect 1146 925 1149 936
rect 1258 933 1276 936
rect 1180 923 1188 926
rect 1260 923 1269 926
rect 1306 925 1309 946
rect 1442 926 1445 936
rect 1508 933 1525 936
rect 1420 925 1445 926
rect 1554 925 1557 936
rect 1594 925 1597 936
rect 1420 923 1444 925
rect 1602 923 1605 934
rect 1690 923 1693 934
rect 1746 926 1749 934
rect 1722 923 1749 926
rect 1802 923 1805 934
rect 1850 926 1853 934
rect 1850 923 1860 926
rect 1300 903 1309 906
rect 14 867 2004 873
rect 1098 816 1101 825
rect 1122 823 1132 826
rect 1146 823 1156 826
rect 1810 816 1813 823
rect 66 813 76 816
rect 122 813 132 816
rect 194 805 197 816
rect 298 813 333 816
rect 426 813 436 816
rect 548 813 557 816
rect 564 813 573 816
rect 612 813 621 816
rect 234 803 242 806
rect 250 803 268 806
rect 330 805 333 813
rect 372 803 389 806
rect 418 803 428 806
rect 618 805 621 813
rect 842 805 845 816
rect 884 813 901 816
rect 986 807 989 816
rect 1034 813 1045 816
rect 1060 813 1084 816
rect 1098 813 1125 816
rect 1188 813 1197 816
rect 1210 813 1221 816
rect 1266 813 1276 816
rect 1314 813 1332 816
rect 1042 807 1045 813
rect 1210 807 1213 813
rect 1068 803 1076 806
rect 1266 805 1269 813
rect 1362 807 1365 816
rect 1402 813 1429 816
rect 1426 807 1429 813
rect 1274 803 1284 806
rect 1300 803 1309 806
rect 1474 805 1477 816
rect 1482 813 1508 816
rect 1570 813 1597 816
rect 1628 813 1645 816
rect 1684 813 1693 816
rect 1716 813 1725 816
rect 1738 813 1748 816
rect 1780 813 1789 816
rect 1810 813 1828 816
rect 1924 813 1941 816
rect 1594 805 1597 813
rect 1650 803 1660 806
rect 1682 803 1692 806
rect 1738 805 1741 813
rect 1746 803 1756 806
rect 1778 803 1788 806
rect 38 767 1980 773
rect 1298 736 1301 745
rect 1506 736 1509 745
rect 1874 736 1877 745
rect 74 723 92 726
rect 186 723 189 734
rect 212 733 221 736
rect 234 726 237 734
rect 282 733 292 736
rect 234 723 245 726
rect 258 723 276 726
rect 314 723 317 734
rect 362 733 372 736
rect 426 723 444 726
rect 578 723 581 734
rect 594 723 597 734
rect 644 723 653 726
rect 722 723 725 734
rect 930 726 933 734
rect 738 723 748 726
rect 914 723 933 726
rect 978 726 981 734
rect 986 733 996 736
rect 1018 733 1028 736
rect 978 723 988 726
rect 1020 723 1029 726
rect 1060 723 1077 726
rect 1082 723 1085 734
rect 1130 726 1133 734
rect 1130 723 1140 726
rect 1170 723 1173 734
rect 1242 723 1245 734
rect 1292 733 1301 736
rect 1322 733 1340 736
rect 1346 733 1364 736
rect 1386 726 1389 736
rect 1268 723 1277 726
rect 1290 723 1300 726
rect 1324 723 1333 726
rect 1386 725 1412 726
rect 1388 723 1412 725
rect 1442 723 1445 734
rect 1500 733 1509 736
rect 1484 723 1509 726
rect 1522 725 1525 736
rect 1580 724 1597 727
rect 1650 726 1653 734
rect 260 713 269 716
rect 1594 715 1597 724
rect 1618 723 1636 726
rect 1642 723 1653 726
rect 1698 723 1701 734
rect 1706 723 1709 734
rect 1754 723 1757 734
rect 1874 733 1892 736
rect 1898 725 1901 736
rect 1932 733 2013 736
rect 1940 723 1949 726
rect 1642 713 1645 723
rect 14 667 2004 673
rect 1252 623 1260 626
rect 1274 623 1284 626
rect 66 613 76 616
rect 210 613 221 616
rect 218 605 221 613
rect 266 603 276 606
rect 290 603 300 606
rect 322 603 340 606
rect 346 603 349 614
rect 500 613 517 616
rect 556 613 565 616
rect 828 613 845 616
rect 1026 613 1044 616
rect 1154 613 1164 616
rect 1186 613 1197 616
rect 1212 613 1236 616
rect 1194 605 1197 613
rect 1220 603 1228 606
rect 1274 603 1277 614
rect 1322 613 1348 616
rect 1450 613 1460 616
rect 1338 605 1341 613
rect 1372 603 1381 606
rect 1450 605 1453 613
rect 1458 603 1468 606
rect 1490 603 1493 614
rect 1548 613 1557 616
rect 1602 613 1628 616
rect 1700 613 1724 616
rect 1796 613 1821 616
rect 1868 613 1885 616
rect 1930 613 2013 616
rect 1540 603 1556 606
rect 1666 603 1676 606
rect 1882 605 1885 613
rect 1932 603 1949 606
rect 38 567 1980 573
rect 538 536 541 545
rect 202 533 212 536
rect 242 526 245 535
rect 284 533 293 536
rect 314 533 324 536
rect 532 533 541 536
rect 650 533 660 536
rect 708 533 717 536
rect 746 533 756 536
rect 836 533 852 536
rect 234 523 245 526
rect 292 523 301 526
rect 322 523 341 526
rect 482 523 485 533
rect 610 526 613 533
rect 610 523 620 526
rect 658 523 676 526
rect 746 525 749 533
rect 906 526 909 533
rect 754 523 780 526
rect 802 523 812 526
rect 898 523 909 526
rect 970 523 973 533
rect 978 523 981 533
rect 1026 523 1060 526
rect 1082 523 1085 533
rect 1106 523 1116 526
rect 1138 525 1141 536
rect 1170 533 1180 536
rect 1306 526 1309 533
rect 1188 523 1197 526
rect 1236 523 1261 526
rect 1290 523 1316 526
rect 1346 525 1349 536
rect 1370 533 1380 536
rect 1506 533 1516 536
rect 1532 533 1548 536
rect 1652 533 1661 536
rect 1372 523 1381 526
rect 1434 523 1437 533
rect 1466 523 1500 526
rect 1540 523 1549 526
rect 1578 523 1620 526
rect 1658 525 1661 533
rect 1690 533 1700 536
rect 1818 533 1828 536
rect 2010 533 2013 613
rect 1690 525 1693 533
rect 1758 523 1765 526
rect 1770 523 1773 533
rect 1826 523 1844 526
rect 1930 523 1933 533
rect 14 467 2004 473
rect 530 453 557 456
rect 530 443 557 446
rect 1322 433 1340 436
rect 1314 423 1324 426
rect 122 413 132 416
rect 266 403 276 406
rect 298 403 308 406
rect 466 405 469 416
rect 490 407 493 416
rect 562 406 565 414
rect 602 413 620 416
rect 658 413 684 416
rect 706 407 709 416
rect 748 413 757 416
rect 530 403 565 406
rect 594 403 604 406
rect 754 405 757 413
rect 802 407 805 416
rect 844 413 853 416
rect 882 413 924 416
rect 1018 414 1036 416
rect 898 407 901 413
rect 836 403 852 406
rect 978 403 988 406
rect 1010 403 1013 414
rect 1018 413 1037 414
rect 1050 413 1060 416
rect 1034 403 1037 413
rect 1074 407 1077 416
rect 1130 413 1141 416
rect 1164 413 1173 416
rect 1130 407 1133 413
rect 1138 407 1141 413
rect 1186 407 1189 416
rect 1228 413 1237 416
rect 1266 413 1292 416
rect 1044 403 1053 406
rect 1194 403 1204 406
rect 1226 403 1236 406
rect 1330 403 1333 414
rect 1354 407 1357 416
rect 1370 413 1380 416
rect 1434 413 1444 416
rect 1404 403 1412 406
rect 1436 403 1445 406
rect 1468 403 1492 406
rect 1514 403 1517 414
rect 1522 405 1525 416
rect 1570 405 1573 416
rect 1578 413 1596 416
rect 1602 405 1605 416
rect 1636 414 1660 416
rect 1636 413 1661 414
rect 1658 403 1661 413
rect 1754 405 1757 416
rect 1762 405 1765 416
rect 1788 414 1820 416
rect 1788 413 1821 414
rect 1818 403 1821 413
rect 1850 403 1853 414
rect 1908 403 1924 406
rect 38 367 1980 373
rect 698 336 701 345
rect 324 333 340 336
rect 346 333 356 336
rect 66 323 92 326
rect 284 323 293 326
rect 348 323 364 326
rect 418 323 428 326
rect 530 323 556 326
rect 586 323 589 334
rect 642 326 645 334
rect 692 333 701 336
rect 708 333 717 336
rect 634 323 645 326
rect 722 323 725 334
rect 778 333 804 336
rect 826 333 836 336
rect 778 326 781 333
rect 748 323 781 326
rect 786 323 796 326
rect 860 323 901 326
rect 906 323 909 334
rect 938 323 980 326
rect 1018 323 1021 334
rect 1212 333 1229 336
rect 1252 333 1277 336
rect 1332 333 1348 336
rect 1372 333 1380 336
rect 1394 333 1420 336
rect 1426 333 1437 336
rect 1466 333 1476 336
rect 1642 333 1652 336
rect 1658 333 1676 336
rect 1690 333 1700 336
rect 1722 333 1732 336
rect 1274 326 1277 333
rect 1130 323 1156 326
rect 1274 323 1300 326
rect 1370 323 1388 326
rect 1426 325 1429 333
rect 1468 323 1477 326
rect 1658 325 1661 333
rect 1690 325 1693 333
rect 1698 323 1708 326
rect 1714 323 1724 326
rect 1754 325 1757 336
rect 1882 326 1885 334
rect 1812 323 1837 326
rect 1882 323 1916 326
rect 1338 313 1348 316
rect 490 303 508 306
rect 14 267 2004 273
rect 540 233 557 236
rect 1010 233 1028 236
rect 1914 233 1924 236
rect 498 216 501 225
rect 522 223 532 226
rect 674 216 677 225
rect 708 223 716 226
rect 1036 223 1044 226
rect 1122 223 1132 226
rect 1698 216 1701 225
rect 74 213 100 216
rect 212 213 221 216
rect 244 213 253 216
rect 276 213 292 216
rect 252 203 268 206
rect 298 203 308 206
rect 330 203 348 206
rect 370 203 373 214
rect 410 203 413 214
rect 418 205 421 216
rect 450 213 469 216
rect 498 213 525 216
rect 466 205 469 213
rect 562 205 565 216
rect 578 213 588 216
rect 610 213 620 216
rect 674 213 692 216
rect 612 203 628 206
rect 674 203 684 206
rect 706 205 709 216
rect 746 213 756 216
rect 810 203 813 214
rect 948 213 957 216
rect 836 203 853 206
rect 954 205 957 213
rect 1042 205 1045 216
rect 1060 213 1077 216
rect 1098 213 1116 216
rect 1186 213 1196 216
rect 1332 213 1341 216
rect 1284 203 1301 206
rect 1386 205 1389 216
rect 1442 205 1445 216
rect 1468 213 1500 216
rect 1530 213 1541 216
rect 1538 205 1541 213
rect 1586 205 1589 216
rect 1642 205 1645 216
rect 1674 213 1692 216
rect 1698 213 1716 216
rect 1676 203 1684 206
rect 1698 203 1708 206
rect 1738 205 1741 216
rect 1786 205 1789 216
rect 1794 205 1797 216
rect 1860 213 1877 216
rect 1866 203 1876 206
rect 38 167 1980 173
rect 274 126 277 134
rect 274 123 284 126
rect 362 123 365 134
rect 466 126 469 134
rect 492 133 501 136
rect 506 133 516 136
rect 396 123 429 126
rect 444 123 460 126
rect 466 123 476 126
rect 530 123 533 134
rect 580 133 596 136
rect 618 133 628 136
rect 546 123 556 126
rect 578 123 588 126
rect 618 125 621 133
rect 626 123 644 126
rect 708 123 733 126
rect 764 123 773 126
rect 818 123 821 134
rect 882 123 885 134
rect 932 133 941 136
rect 964 134 980 136
rect 964 133 981 134
rect 1028 133 1037 136
rect 938 125 941 133
rect 978 123 981 133
rect 1004 123 1029 126
rect 1068 123 1092 126
rect 1122 123 1125 134
rect 1130 123 1133 134
rect 1226 126 1229 134
rect 1164 123 1181 126
rect 1220 123 1229 126
rect 1322 123 1325 134
rect 1372 133 1380 136
rect 1492 133 1500 136
rect 1522 123 1525 134
rect 1530 123 1540 126
rect 1554 123 1557 134
rect 1610 123 1613 134
rect 1818 133 1828 136
rect 1852 133 1860 136
rect 1642 123 1668 126
rect 1730 123 1756 126
rect 1820 123 1829 126
rect 1906 123 1909 134
rect 1690 113 1700 116
rect 1410 103 1428 106
rect 1690 103 1716 106
rect 14 67 2004 73
rect 38 37 1980 57
rect 14 13 2004 33
<< metal2 >>
rect 14 13 34 1927
rect 38 37 58 1903
rect 74 1813 85 1816
rect 130 1793 133 1816
rect 66 1723 69 1736
rect 130 1723 133 1746
rect 66 1533 69 1616
rect 130 1613 133 1626
rect 66 1293 69 1526
rect 82 1426 85 1526
rect 82 1423 93 1426
rect 74 1333 77 1416
rect 90 1356 93 1423
rect 130 1413 133 1526
rect 154 1523 157 1806
rect 170 1803 173 1816
rect 178 1813 181 1836
rect 210 1823 213 1836
rect 234 1833 253 1836
rect 202 1756 205 1806
rect 210 1793 213 1806
rect 226 1756 229 1816
rect 234 1803 237 1833
rect 202 1753 213 1756
rect 226 1753 237 1756
rect 170 1733 181 1736
rect 186 1733 189 1746
rect 210 1726 213 1753
rect 186 1723 205 1726
rect 210 1723 221 1726
rect 234 1723 237 1753
rect 186 1703 189 1716
rect 218 1713 221 1723
rect 170 1613 173 1626
rect 178 1603 181 1616
rect 186 1566 189 1616
rect 226 1613 229 1706
rect 234 1703 237 1716
rect 242 1713 245 1826
rect 250 1653 253 1833
rect 322 1833 333 1836
rect 322 1826 325 1833
rect 266 1816 269 1826
rect 258 1803 261 1816
rect 266 1813 277 1816
rect 290 1813 293 1826
rect 306 1823 325 1826
rect 258 1723 269 1726
rect 266 1713 269 1723
rect 274 1666 277 1806
rect 282 1676 285 1806
rect 298 1743 301 1816
rect 306 1803 309 1816
rect 322 1773 325 1823
rect 298 1723 301 1736
rect 306 1733 309 1766
rect 330 1763 333 1826
rect 338 1813 341 1826
rect 290 1693 293 1716
rect 322 1713 325 1726
rect 282 1673 301 1676
rect 274 1663 293 1666
rect 242 1613 253 1616
rect 266 1593 269 1636
rect 282 1623 285 1656
rect 290 1613 293 1663
rect 298 1633 301 1673
rect 338 1633 341 1734
rect 354 1703 357 1826
rect 362 1793 365 1816
rect 386 1746 389 1766
rect 402 1753 405 1816
rect 442 1786 445 1806
rect 466 1786 469 1806
rect 442 1783 469 1786
rect 442 1763 445 1783
rect 378 1743 389 1746
rect 362 1646 365 1726
rect 378 1686 381 1743
rect 378 1683 389 1686
rect 354 1643 365 1646
rect 306 1623 349 1626
rect 306 1613 317 1616
rect 330 1613 333 1623
rect 322 1603 333 1606
rect 186 1563 197 1566
rect 178 1436 181 1536
rect 194 1473 197 1563
rect 218 1513 221 1526
rect 162 1433 181 1436
rect 138 1376 141 1416
rect 138 1373 149 1376
rect 82 1353 93 1356
rect 66 1213 69 1226
rect 82 1183 85 1353
rect 90 1313 93 1326
rect 98 1276 101 1336
rect 114 1326 117 1366
rect 106 1323 117 1326
rect 122 1323 125 1356
rect 130 1326 133 1336
rect 146 1333 149 1373
rect 162 1356 165 1433
rect 154 1353 165 1356
rect 130 1323 149 1326
rect 114 1286 117 1323
rect 114 1283 125 1286
rect 98 1273 117 1276
rect 114 1213 117 1273
rect 114 1166 117 1186
rect 110 1163 117 1166
rect 66 1013 69 1156
rect 74 1073 77 1126
rect 110 1116 113 1163
rect 122 1123 125 1283
rect 130 1223 133 1323
rect 154 1256 157 1353
rect 162 1343 173 1346
rect 162 1263 165 1316
rect 170 1303 173 1326
rect 138 1253 157 1256
rect 138 1176 141 1253
rect 154 1183 157 1206
rect 138 1173 157 1176
rect 130 1123 133 1146
rect 110 1113 117 1116
rect 74 983 77 1036
rect 114 1013 117 1113
rect 154 1096 157 1173
rect 170 1156 173 1226
rect 178 1216 181 1406
rect 186 1223 189 1336
rect 194 1333 197 1416
rect 202 1363 205 1486
rect 218 1423 221 1456
rect 218 1403 221 1416
rect 258 1413 261 1546
rect 282 1543 293 1546
rect 274 1453 277 1526
rect 282 1483 285 1526
rect 290 1513 293 1536
rect 282 1413 285 1476
rect 306 1446 309 1546
rect 314 1473 317 1526
rect 322 1523 325 1536
rect 338 1533 341 1546
rect 346 1533 349 1616
rect 354 1613 357 1643
rect 330 1523 341 1526
rect 338 1493 341 1516
rect 298 1443 309 1446
rect 202 1333 205 1346
rect 226 1326 229 1406
rect 274 1346 277 1406
rect 250 1343 277 1346
rect 194 1216 197 1236
rect 202 1226 205 1326
rect 210 1283 213 1326
rect 218 1323 229 1326
rect 202 1223 213 1226
rect 178 1213 189 1216
rect 194 1213 205 1216
rect 170 1153 181 1156
rect 170 1133 173 1146
rect 178 1126 181 1153
rect 194 1133 197 1206
rect 202 1203 205 1213
rect 210 1196 213 1223
rect 218 1213 221 1323
rect 226 1203 229 1316
rect 170 1123 181 1126
rect 170 1113 173 1123
rect 154 1093 181 1096
rect 130 993 133 1016
rect 74 913 77 956
rect 66 813 69 856
rect 66 696 69 756
rect 74 723 77 876
rect 122 813 125 946
rect 130 923 133 936
rect 138 883 141 966
rect 154 953 157 1016
rect 170 1003 173 1076
rect 154 856 157 936
rect 170 933 173 946
rect 170 903 173 916
rect 138 853 157 856
rect 138 836 141 853
rect 178 846 181 1093
rect 186 1016 189 1126
rect 202 1053 205 1196
rect 210 1193 229 1196
rect 226 1183 229 1193
rect 234 1176 237 1286
rect 242 1213 245 1326
rect 250 1293 253 1343
rect 282 1333 285 1346
rect 290 1333 293 1416
rect 298 1343 301 1443
rect 306 1423 309 1436
rect 314 1413 325 1416
rect 306 1403 333 1406
rect 338 1383 341 1446
rect 346 1403 349 1526
rect 354 1413 357 1516
rect 362 1513 365 1616
rect 386 1553 389 1683
rect 402 1613 405 1716
rect 418 1693 421 1736
rect 426 1633 429 1746
rect 474 1733 477 1776
rect 482 1733 485 1746
rect 490 1733 493 1940
rect 522 1856 525 1940
rect 570 1926 573 1940
rect 514 1853 525 1856
rect 562 1923 573 1926
rect 506 1803 509 1816
rect 514 1793 517 1853
rect 506 1726 509 1736
rect 514 1733 517 1746
rect 530 1733 533 1806
rect 546 1803 549 1816
rect 554 1793 557 1806
rect 562 1773 565 1923
rect 586 1856 589 1940
rect 602 1926 605 1940
rect 602 1923 613 1926
rect 586 1853 597 1856
rect 570 1813 581 1816
rect 546 1726 549 1736
rect 554 1733 557 1746
rect 482 1723 509 1726
rect 370 1423 373 1526
rect 378 1446 381 1536
rect 386 1523 397 1526
rect 394 1503 397 1516
rect 402 1513 405 1526
rect 410 1523 413 1616
rect 418 1526 421 1626
rect 450 1606 453 1706
rect 482 1703 485 1716
rect 514 1713 517 1726
rect 522 1703 525 1726
rect 530 1723 541 1726
rect 546 1723 557 1726
rect 562 1696 565 1756
rect 570 1703 573 1796
rect 578 1733 581 1806
rect 586 1793 589 1806
rect 594 1803 597 1853
rect 610 1836 613 1923
rect 658 1856 661 1940
rect 650 1853 661 1856
rect 610 1833 621 1836
rect 602 1803 605 1816
rect 610 1813 613 1826
rect 610 1793 613 1806
rect 618 1786 621 1833
rect 602 1783 621 1786
rect 578 1713 581 1726
rect 530 1656 533 1696
rect 562 1693 573 1696
rect 522 1653 533 1656
rect 434 1603 453 1606
rect 426 1533 429 1546
rect 418 1523 429 1526
rect 426 1513 429 1523
rect 378 1443 397 1446
rect 442 1443 445 1596
rect 458 1573 461 1616
rect 466 1613 469 1626
rect 482 1583 485 1616
rect 506 1613 509 1626
rect 522 1576 525 1653
rect 522 1573 533 1576
rect 466 1523 469 1546
rect 482 1536 485 1556
rect 482 1533 489 1536
rect 530 1533 533 1573
rect 258 1286 261 1326
rect 274 1313 277 1326
rect 282 1313 285 1326
rect 290 1323 301 1326
rect 306 1306 309 1326
rect 322 1323 333 1326
rect 322 1313 333 1316
rect 266 1303 277 1306
rect 306 1303 317 1306
rect 250 1283 261 1286
rect 250 1213 253 1283
rect 210 1046 213 1136
rect 218 1103 221 1176
rect 226 1173 237 1176
rect 226 1153 229 1173
rect 242 1166 245 1206
rect 234 1163 245 1166
rect 234 1136 237 1163
rect 230 1133 237 1136
rect 250 1136 253 1206
rect 266 1193 269 1296
rect 274 1283 277 1303
rect 274 1183 277 1196
rect 282 1173 285 1206
rect 290 1196 293 1236
rect 298 1213 301 1226
rect 306 1203 309 1236
rect 314 1203 317 1216
rect 290 1193 317 1196
rect 322 1143 325 1296
rect 338 1266 341 1316
rect 346 1273 349 1326
rect 338 1263 349 1266
rect 250 1133 261 1136
rect 230 1086 233 1133
rect 258 1086 261 1133
rect 274 1113 277 1126
rect 298 1093 301 1136
rect 314 1113 317 1136
rect 322 1113 325 1126
rect 230 1083 237 1086
rect 210 1043 221 1046
rect 186 1013 213 1016
rect 186 993 189 1006
rect 218 1003 221 1043
rect 234 1026 237 1083
rect 250 1083 261 1086
rect 226 993 229 1026
rect 234 1023 245 1026
rect 194 933 197 946
rect 134 833 141 836
rect 154 843 181 846
rect 134 746 137 833
rect 134 743 141 746
rect 130 706 133 726
rect 138 713 141 743
rect 146 723 149 746
rect 154 706 157 843
rect 170 816 173 826
rect 170 813 181 816
rect 170 743 173 806
rect 178 803 181 813
rect 186 796 189 926
rect 194 903 197 926
rect 202 853 205 916
rect 194 813 197 826
rect 202 813 205 826
rect 194 803 205 806
rect 186 793 205 796
rect 126 703 133 706
rect 138 703 157 706
rect 66 693 85 696
rect 66 613 69 686
rect 82 606 85 693
rect 74 603 85 606
rect 74 503 77 603
rect 106 513 109 676
rect 126 636 129 703
rect 126 633 133 636
rect 114 473 117 626
rect 130 613 133 633
rect 138 576 141 703
rect 170 636 173 736
rect 186 723 197 726
rect 186 643 189 716
rect 154 633 173 636
rect 154 603 157 633
rect 186 616 189 626
rect 138 573 157 576
rect 74 463 85 466
rect 74 413 77 463
rect 122 413 125 536
rect 130 524 133 566
rect 138 456 141 546
rect 134 453 141 456
rect 154 453 157 573
rect 170 533 173 616
rect 186 613 197 616
rect 202 613 205 793
rect 210 773 213 986
rect 226 933 229 966
rect 234 933 237 1016
rect 242 946 245 1023
rect 250 1003 253 1083
rect 330 1076 333 1226
rect 338 1183 341 1256
rect 346 1223 349 1263
rect 346 1203 349 1216
rect 354 1213 357 1326
rect 362 1293 365 1416
rect 370 1366 373 1416
rect 378 1413 381 1436
rect 386 1406 389 1426
rect 378 1403 389 1406
rect 394 1403 397 1443
rect 418 1423 437 1426
rect 370 1363 381 1366
rect 362 1206 365 1276
rect 378 1253 381 1363
rect 386 1263 389 1296
rect 378 1213 381 1246
rect 362 1203 381 1206
rect 314 1073 333 1076
rect 258 1023 269 1026
rect 258 1013 261 1023
rect 266 996 269 1016
rect 274 1013 277 1036
rect 266 993 277 996
rect 242 943 261 946
rect 242 933 253 936
rect 218 766 221 926
rect 242 916 245 926
rect 226 913 245 916
rect 250 913 253 926
rect 226 833 229 913
rect 258 906 261 943
rect 242 903 261 906
rect 226 783 229 806
rect 234 803 237 886
rect 234 773 237 796
rect 218 763 237 766
rect 218 733 229 736
rect 218 713 221 726
rect 210 613 213 646
rect 218 613 221 686
rect 178 546 181 606
rect 186 563 189 606
rect 194 576 197 613
rect 210 583 213 606
rect 194 573 205 576
rect 178 543 189 546
rect 170 493 173 526
rect 74 366 77 386
rect 134 376 137 453
rect 154 403 157 426
rect 178 413 181 536
rect 186 523 189 543
rect 194 463 197 536
rect 202 533 205 573
rect 210 573 221 576
rect 178 386 181 406
rect 194 393 197 456
rect 202 426 205 526
rect 210 503 213 573
rect 226 556 229 726
rect 234 706 237 763
rect 242 723 245 903
rect 266 893 269 976
rect 274 933 277 993
rect 282 933 285 1006
rect 290 1003 293 1016
rect 298 1013 301 1056
rect 298 993 301 1006
rect 282 923 293 926
rect 274 913 285 916
rect 298 903 301 926
rect 250 816 253 836
rect 250 813 269 816
rect 250 783 253 806
rect 258 773 261 796
rect 266 763 269 813
rect 274 803 277 816
rect 234 703 241 706
rect 238 636 241 703
rect 234 633 241 636
rect 234 566 237 633
rect 242 593 245 606
rect 250 603 253 736
rect 258 623 261 726
rect 266 713 269 746
rect 274 706 277 776
rect 282 723 285 896
rect 266 703 277 706
rect 282 703 285 716
rect 266 663 269 703
rect 290 676 293 816
rect 298 813 301 826
rect 298 793 301 806
rect 306 743 309 1006
rect 314 993 317 1073
rect 338 1053 341 1146
rect 346 1113 349 1136
rect 354 1123 357 1136
rect 354 1046 357 1116
rect 322 993 325 1006
rect 330 1003 333 1016
rect 314 943 317 986
rect 338 983 341 1016
rect 314 893 317 936
rect 330 933 333 946
rect 330 856 333 926
rect 346 903 349 1046
rect 354 1043 365 1046
rect 370 1043 373 1186
rect 378 1133 381 1196
rect 386 1156 389 1236
rect 394 1203 397 1326
rect 402 1253 405 1416
rect 418 1413 421 1423
rect 410 1403 421 1406
rect 426 1393 429 1416
rect 434 1413 437 1423
rect 434 1403 445 1406
rect 450 1403 453 1416
rect 458 1413 461 1446
rect 402 1223 405 1246
rect 386 1153 397 1156
rect 386 1133 389 1146
rect 354 876 357 1036
rect 362 1003 365 1043
rect 386 1016 389 1066
rect 394 1043 397 1153
rect 402 1123 405 1206
rect 410 1196 413 1316
rect 426 1313 429 1386
rect 418 1203 421 1266
rect 426 1213 429 1286
rect 410 1193 429 1196
rect 426 1176 429 1193
rect 434 1183 437 1206
rect 442 1193 445 1326
rect 458 1323 461 1406
rect 466 1393 469 1406
rect 474 1403 477 1516
rect 486 1436 489 1533
rect 522 1493 525 1526
rect 482 1433 489 1436
rect 482 1403 485 1433
rect 522 1423 525 1436
rect 530 1423 533 1526
rect 538 1416 541 1436
rect 490 1366 493 1416
rect 506 1413 525 1416
rect 530 1413 541 1416
rect 546 1413 549 1516
rect 554 1513 557 1536
rect 562 1503 565 1686
rect 570 1613 573 1693
rect 586 1683 589 1776
rect 602 1733 605 1783
rect 610 1743 613 1756
rect 610 1693 613 1736
rect 618 1733 621 1746
rect 626 1733 629 1816
rect 650 1813 653 1853
rect 658 1813 661 1836
rect 666 1833 685 1836
rect 666 1806 669 1833
rect 642 1793 645 1806
rect 650 1803 669 1806
rect 674 1803 677 1826
rect 682 1803 685 1833
rect 690 1816 693 1836
rect 730 1816 733 1846
rect 690 1813 701 1816
rect 642 1733 645 1756
rect 650 1726 653 1803
rect 682 1783 685 1796
rect 698 1766 701 1813
rect 690 1763 701 1766
rect 626 1723 653 1726
rect 642 1703 645 1716
rect 650 1713 653 1723
rect 658 1716 661 1736
rect 666 1723 669 1746
rect 682 1743 685 1756
rect 658 1713 669 1716
rect 674 1713 677 1736
rect 682 1713 685 1726
rect 666 1706 669 1713
rect 658 1693 661 1706
rect 666 1703 685 1706
rect 690 1703 693 1763
rect 714 1746 717 1816
rect 698 1733 701 1746
rect 706 1743 717 1746
rect 722 1813 733 1816
rect 722 1743 725 1813
rect 706 1723 709 1743
rect 626 1613 629 1626
rect 650 1566 653 1606
rect 650 1563 661 1566
rect 578 1533 581 1546
rect 570 1433 573 1526
rect 594 1456 597 1536
rect 618 1513 621 1526
rect 590 1453 597 1456
rect 562 1423 573 1426
rect 498 1393 501 1406
rect 530 1403 533 1413
rect 546 1393 549 1406
rect 490 1363 501 1366
rect 474 1336 477 1356
rect 474 1333 481 1336
rect 458 1303 461 1316
rect 466 1263 469 1326
rect 478 1266 481 1333
rect 498 1286 501 1363
rect 546 1333 549 1376
rect 554 1353 557 1406
rect 562 1343 565 1423
rect 570 1363 573 1416
rect 578 1346 581 1416
rect 590 1396 593 1453
rect 590 1393 597 1396
rect 594 1373 597 1393
rect 578 1343 589 1346
rect 474 1263 481 1266
rect 490 1283 501 1286
rect 410 1133 413 1146
rect 410 1113 413 1126
rect 418 1116 421 1176
rect 426 1173 445 1176
rect 426 1123 429 1136
rect 418 1113 429 1116
rect 370 993 373 1016
rect 378 1013 389 1016
rect 378 983 381 1013
rect 386 993 389 1006
rect 370 943 389 946
rect 362 913 365 936
rect 370 923 373 943
rect 378 923 381 936
rect 386 933 389 943
rect 394 926 397 986
rect 402 933 405 1006
rect 418 973 421 1056
rect 426 1026 429 1113
rect 434 1033 437 1136
rect 426 1023 437 1026
rect 426 1003 429 1016
rect 386 923 397 926
rect 314 853 333 856
rect 346 873 357 876
rect 314 733 317 853
rect 322 793 325 846
rect 274 673 293 676
rect 258 613 269 616
rect 234 563 245 566
rect 218 553 229 556
rect 218 516 221 553
rect 226 523 229 546
rect 234 534 237 556
rect 242 543 245 563
rect 258 536 261 613
rect 266 593 269 606
rect 274 583 277 673
rect 282 576 285 666
rect 290 613 293 646
rect 298 613 301 726
rect 306 713 309 726
rect 314 696 317 726
rect 306 693 317 696
rect 306 613 309 693
rect 314 616 317 666
rect 322 623 325 726
rect 314 613 325 616
rect 274 573 285 576
rect 290 573 293 606
rect 274 563 277 573
rect 298 566 301 606
rect 314 593 317 606
rect 282 563 301 566
rect 242 533 261 536
rect 266 534 269 546
rect 234 516 237 526
rect 218 513 237 516
rect 226 483 229 506
rect 202 423 213 426
rect 170 383 181 386
rect 134 373 141 376
rect 66 323 69 366
rect 74 363 85 366
rect 82 256 85 363
rect 138 353 141 373
rect 146 323 149 346
rect 170 276 173 383
rect 202 333 205 416
rect 210 383 213 423
rect 202 313 205 326
rect 170 273 181 276
rect 74 253 85 256
rect 74 213 77 253
rect 154 193 157 216
rect 178 203 181 273
rect 194 213 197 226
rect 218 213 221 476
rect 234 466 237 513
rect 242 496 245 533
rect 250 513 253 526
rect 258 496 261 526
rect 274 523 277 536
rect 282 516 285 563
rect 306 556 309 566
rect 298 553 309 556
rect 278 513 285 516
rect 242 493 249 496
rect 258 493 269 496
rect 226 463 237 466
rect 226 333 229 463
rect 246 426 249 493
rect 242 423 249 426
rect 242 373 245 423
rect 258 406 261 486
rect 266 413 269 493
rect 278 436 281 513
rect 290 503 293 536
rect 274 433 281 436
rect 250 403 261 406
rect 250 366 253 403
rect 242 363 253 366
rect 234 323 237 336
rect 242 316 245 363
rect 234 313 245 316
rect 250 296 253 356
rect 258 333 261 396
rect 266 363 269 406
rect 274 386 277 433
rect 282 396 285 416
rect 290 403 293 436
rect 298 413 301 553
rect 298 396 301 406
rect 282 393 301 396
rect 306 393 309 536
rect 314 533 317 586
rect 322 553 325 606
rect 330 603 333 826
rect 338 743 341 816
rect 346 813 349 873
rect 354 803 357 816
rect 362 803 365 816
rect 346 743 365 746
rect 338 683 341 736
rect 346 723 349 743
rect 354 703 357 736
rect 362 733 365 743
rect 362 676 365 726
rect 370 723 373 886
rect 386 876 389 923
rect 402 913 405 926
rect 418 903 421 956
rect 434 883 437 1023
rect 442 953 445 1173
rect 450 983 453 1226
rect 458 1193 461 1206
rect 458 1123 461 1176
rect 466 1133 469 1206
rect 474 1133 477 1263
rect 482 1213 485 1246
rect 490 1176 493 1283
rect 498 1213 501 1266
rect 482 1173 493 1176
rect 482 1133 485 1146
rect 458 1103 461 1116
rect 482 1113 485 1126
rect 490 1073 493 1126
rect 498 1113 501 1166
rect 506 1123 509 1226
rect 514 1213 517 1326
rect 530 1213 533 1226
rect 538 1213 541 1286
rect 546 1223 549 1326
rect 522 1143 525 1206
rect 530 1136 533 1186
rect 546 1183 549 1216
rect 554 1163 557 1256
rect 562 1223 565 1336
rect 570 1303 573 1326
rect 578 1323 581 1336
rect 586 1316 589 1343
rect 578 1313 589 1316
rect 578 1266 581 1313
rect 594 1273 597 1356
rect 602 1333 605 1346
rect 610 1313 613 1336
rect 618 1293 621 1386
rect 578 1263 589 1266
rect 530 1133 549 1136
rect 562 1133 565 1216
rect 578 1166 581 1206
rect 586 1203 589 1263
rect 594 1196 597 1216
rect 602 1203 605 1236
rect 610 1196 613 1206
rect 594 1193 613 1196
rect 618 1166 621 1216
rect 626 1206 629 1506
rect 658 1496 661 1563
rect 666 1543 669 1616
rect 674 1613 677 1626
rect 682 1623 685 1703
rect 674 1523 677 1606
rect 698 1603 701 1626
rect 714 1613 717 1736
rect 722 1693 725 1736
rect 730 1713 733 1806
rect 738 1783 741 1836
rect 754 1823 757 1836
rect 738 1703 741 1726
rect 746 1703 749 1816
rect 754 1793 757 1806
rect 754 1713 757 1786
rect 762 1766 765 1876
rect 770 1806 773 1856
rect 786 1823 789 1836
rect 802 1823 805 1836
rect 810 1823 813 1856
rect 778 1813 821 1816
rect 770 1803 781 1806
rect 762 1763 773 1766
rect 762 1733 765 1756
rect 762 1713 765 1726
rect 770 1716 773 1763
rect 778 1726 781 1803
rect 786 1733 789 1746
rect 778 1723 789 1726
rect 770 1713 781 1716
rect 786 1713 789 1723
rect 778 1656 781 1713
rect 778 1653 785 1656
rect 714 1583 717 1606
rect 730 1583 733 1646
rect 738 1616 741 1636
rect 738 1613 749 1616
rect 682 1533 685 1546
rect 714 1533 717 1546
rect 722 1543 733 1546
rect 682 1503 685 1526
rect 634 1333 637 1416
rect 634 1313 637 1326
rect 642 1263 645 1496
rect 658 1493 685 1496
rect 722 1493 725 1543
rect 730 1513 733 1536
rect 738 1523 741 1606
rect 746 1543 749 1613
rect 782 1596 785 1653
rect 794 1613 797 1776
rect 802 1633 805 1806
rect 826 1773 829 1940
rect 842 1873 845 1940
rect 858 1836 861 1940
rect 834 1823 837 1836
rect 850 1833 861 1836
rect 850 1826 853 1833
rect 842 1823 853 1826
rect 810 1733 813 1756
rect 834 1753 837 1806
rect 842 1786 845 1823
rect 850 1793 853 1816
rect 858 1803 861 1826
rect 866 1816 869 1856
rect 874 1823 877 1940
rect 890 1826 893 1940
rect 906 1873 909 1940
rect 898 1833 901 1866
rect 922 1863 925 1940
rect 938 1883 941 1940
rect 954 1893 957 1940
rect 970 1903 973 1940
rect 890 1823 909 1826
rect 866 1813 901 1816
rect 842 1783 861 1786
rect 834 1723 837 1746
rect 858 1743 861 1783
rect 866 1773 869 1796
rect 858 1723 861 1736
rect 866 1733 877 1736
rect 882 1733 885 1806
rect 890 1743 893 1813
rect 906 1733 909 1823
rect 914 1813 917 1826
rect 922 1803 925 1826
rect 930 1813 933 1846
rect 938 1816 941 1826
rect 938 1813 949 1816
rect 954 1813 957 1836
rect 938 1793 941 1806
rect 946 1796 949 1813
rect 962 1803 965 1826
rect 970 1803 973 1846
rect 978 1813 981 1826
rect 994 1816 997 1826
rect 986 1813 997 1816
rect 946 1793 965 1796
rect 938 1743 941 1756
rect 802 1613 805 1626
rect 834 1613 837 1626
rect 778 1593 785 1596
rect 778 1576 781 1593
rect 802 1583 805 1596
rect 770 1573 781 1576
rect 650 1333 653 1346
rect 658 1333 661 1436
rect 682 1343 685 1493
rect 770 1486 773 1573
rect 818 1553 821 1606
rect 842 1596 845 1616
rect 850 1613 853 1636
rect 858 1603 861 1716
rect 866 1613 869 1733
rect 874 1696 877 1726
rect 882 1713 885 1726
rect 914 1723 917 1736
rect 874 1693 885 1696
rect 842 1593 869 1596
rect 882 1586 885 1693
rect 898 1613 901 1636
rect 914 1623 941 1626
rect 874 1583 885 1586
rect 898 1583 901 1606
rect 778 1513 781 1526
rect 762 1483 773 1486
rect 666 1333 685 1336
rect 658 1263 661 1326
rect 666 1283 669 1333
rect 674 1256 677 1326
rect 682 1313 685 1326
rect 690 1293 693 1326
rect 658 1236 661 1256
rect 674 1253 685 1256
rect 634 1213 637 1226
rect 626 1203 637 1206
rect 578 1163 585 1166
rect 522 1103 525 1126
rect 530 1113 533 1126
rect 466 1026 469 1046
rect 466 1023 477 1026
rect 474 976 477 1023
rect 490 993 493 1006
rect 498 1003 501 1016
rect 466 973 477 976
rect 514 976 517 1096
rect 546 1093 549 1126
rect 582 1106 585 1163
rect 578 1103 585 1106
rect 594 1163 621 1166
rect 514 973 533 976
rect 466 946 469 973
rect 458 943 469 946
rect 458 926 461 943
rect 442 913 445 926
rect 454 923 461 926
rect 378 873 389 876
rect 378 736 381 873
rect 454 866 457 923
rect 454 863 461 866
rect 386 813 389 826
rect 386 783 389 806
rect 394 803 397 856
rect 458 843 461 863
rect 402 796 405 816
rect 410 803 413 816
rect 418 813 421 836
rect 418 796 421 806
rect 402 793 421 796
rect 426 773 429 816
rect 450 813 453 826
rect 434 803 445 806
rect 466 776 469 936
rect 490 923 501 926
rect 514 923 517 936
rect 482 806 485 906
rect 530 856 533 973
rect 546 966 549 1036
rect 554 993 557 1016
rect 546 963 557 966
rect 554 886 557 963
rect 570 923 573 946
rect 546 883 557 886
rect 490 813 493 826
rect 482 803 493 806
rect 450 773 469 776
rect 378 733 397 736
rect 378 713 381 726
rect 386 703 389 726
rect 394 693 397 733
rect 346 673 365 676
rect 346 646 349 673
rect 338 643 349 646
rect 338 596 341 643
rect 330 593 341 596
rect 346 546 349 606
rect 322 543 349 546
rect 314 456 317 526
rect 322 523 325 543
rect 330 533 341 536
rect 330 463 333 526
rect 338 483 341 526
rect 346 513 349 526
rect 314 453 325 456
rect 314 413 317 426
rect 330 403 333 416
rect 354 413 357 426
rect 362 413 365 666
rect 378 486 381 616
rect 386 613 389 626
rect 386 513 389 526
rect 394 493 397 606
rect 402 486 405 736
rect 426 713 429 726
rect 370 483 381 486
rect 394 483 405 486
rect 274 383 281 386
rect 266 333 269 346
rect 266 313 269 326
rect 278 296 281 383
rect 290 333 293 346
rect 290 303 293 326
rect 298 323 301 336
rect 306 316 309 366
rect 298 313 309 316
rect 314 313 317 326
rect 242 293 253 296
rect 242 236 245 293
rect 226 223 229 236
rect 242 233 253 236
rect 194 193 197 206
rect 218 183 221 206
rect 226 203 229 216
rect 250 213 253 233
rect 226 133 229 196
rect 258 193 261 296
rect 278 293 285 296
rect 258 113 261 126
rect 274 113 277 216
rect 282 183 285 293
rect 290 206 293 226
rect 298 213 309 216
rect 314 213 317 246
rect 290 203 301 206
rect 290 113 293 156
rect 314 146 317 206
rect 322 183 325 376
rect 330 293 333 386
rect 346 333 349 346
rect 330 213 333 286
rect 338 213 341 226
rect 330 153 333 206
rect 346 153 349 326
rect 354 313 357 406
rect 370 343 373 483
rect 378 403 381 446
rect 394 383 397 483
rect 402 363 405 426
rect 410 413 413 556
rect 426 486 429 676
rect 418 483 429 486
rect 418 413 421 483
rect 434 473 437 766
rect 442 593 445 696
rect 450 663 453 773
rect 490 756 493 803
rect 466 753 493 756
rect 466 733 469 753
rect 490 733 493 753
rect 458 613 461 626
rect 450 553 453 606
rect 474 603 477 656
rect 506 626 509 856
rect 530 853 537 856
rect 514 723 517 776
rect 534 766 537 853
rect 502 623 509 626
rect 458 583 469 586
rect 442 513 445 546
rect 450 523 453 536
rect 458 523 461 583
rect 502 576 505 623
rect 514 593 517 616
rect 522 613 525 766
rect 530 763 537 766
rect 546 763 549 883
rect 578 833 581 1103
rect 586 996 589 1086
rect 594 1063 597 1163
rect 602 1123 605 1146
rect 594 1013 597 1036
rect 594 1003 605 1006
rect 586 993 601 996
rect 598 856 601 993
rect 610 986 613 1156
rect 642 1153 645 1216
rect 650 1133 653 1236
rect 658 1233 665 1236
rect 642 1083 645 1126
rect 618 993 621 1006
rect 626 1003 629 1016
rect 642 1013 645 1066
rect 650 1006 653 1126
rect 662 1066 665 1233
rect 682 1213 685 1253
rect 690 1213 693 1226
rect 674 1123 677 1156
rect 682 1133 685 1146
rect 698 1143 701 1446
rect 706 1333 709 1416
rect 714 1343 717 1386
rect 706 1313 709 1326
rect 706 1193 709 1226
rect 714 1176 717 1296
rect 722 1253 725 1346
rect 730 1293 733 1326
rect 738 1286 741 1376
rect 746 1323 749 1356
rect 762 1346 765 1483
rect 818 1466 821 1536
rect 834 1523 837 1546
rect 874 1523 877 1583
rect 906 1563 909 1616
rect 914 1613 917 1623
rect 922 1576 925 1616
rect 930 1583 933 1606
rect 914 1573 925 1576
rect 826 1486 829 1506
rect 826 1483 837 1486
rect 810 1463 821 1466
rect 754 1343 765 1346
rect 770 1346 773 1396
rect 786 1393 789 1416
rect 770 1343 781 1346
rect 754 1316 757 1343
rect 762 1323 765 1336
rect 754 1313 765 1316
rect 730 1283 741 1286
rect 730 1203 733 1283
rect 762 1273 765 1313
rect 754 1203 757 1216
rect 714 1173 733 1176
rect 690 1106 693 1126
rect 698 1123 701 1136
rect 706 1133 725 1136
rect 706 1113 709 1133
rect 634 1003 653 1006
rect 610 983 629 986
rect 610 933 621 936
rect 598 853 605 856
rect 554 783 557 816
rect 570 813 573 826
rect 578 813 589 816
rect 594 813 597 836
rect 562 803 573 806
rect 586 803 597 806
rect 530 653 533 763
rect 502 573 509 576
rect 466 533 469 546
rect 466 516 469 526
rect 474 523 477 566
rect 506 556 509 573
rect 498 553 509 556
rect 530 533 533 546
rect 466 513 477 516
rect 482 513 485 526
rect 442 443 445 496
rect 442 413 445 426
rect 450 413 453 506
rect 466 413 469 466
rect 474 443 477 513
rect 498 503 501 526
rect 514 436 517 526
rect 522 453 533 456
rect 522 443 525 453
rect 410 386 413 406
rect 418 393 421 406
rect 410 383 437 386
rect 370 303 373 336
rect 418 333 421 346
rect 386 283 389 326
rect 402 276 405 326
rect 418 303 421 326
rect 426 323 429 366
rect 354 213 357 276
rect 402 273 409 276
rect 362 203 365 216
rect 378 213 381 226
rect 394 213 397 266
rect 406 226 409 273
rect 434 253 437 383
rect 442 236 445 326
rect 402 223 409 226
rect 418 233 445 236
rect 370 183 373 206
rect 386 163 389 206
rect 402 203 405 223
rect 418 213 421 233
rect 442 213 445 226
rect 450 213 453 336
rect 458 333 461 346
rect 458 303 461 316
rect 458 263 461 286
rect 410 183 413 206
rect 298 143 317 146
rect 298 123 301 143
rect 306 103 309 136
rect 314 133 317 143
rect 370 133 373 146
rect 338 113 341 126
rect 362 103 365 126
rect 418 123 421 136
rect 426 133 429 146
rect 434 126 437 166
rect 450 133 453 166
rect 426 123 437 126
rect 458 123 461 186
rect 466 173 469 406
rect 474 323 477 436
rect 506 433 517 436
rect 482 386 485 416
rect 490 413 493 426
rect 498 416 501 426
rect 498 413 509 416
rect 514 413 517 433
rect 506 406 509 413
rect 498 393 501 406
rect 506 403 517 406
rect 482 383 501 386
rect 482 333 485 346
rect 490 313 493 366
rect 490 293 493 306
rect 498 303 501 383
rect 506 306 509 386
rect 514 313 517 403
rect 522 343 525 426
rect 530 413 533 446
rect 530 333 533 406
rect 538 373 541 746
rect 554 676 557 776
rect 550 673 557 676
rect 562 673 565 796
rect 570 723 573 803
rect 602 773 605 853
rect 610 793 613 926
rect 618 763 621 926
rect 626 916 629 983
rect 634 933 637 946
rect 642 926 645 996
rect 634 923 645 926
rect 626 913 645 916
rect 626 766 629 906
rect 634 803 637 816
rect 626 763 637 766
rect 578 713 581 726
rect 586 723 589 756
rect 594 693 597 726
rect 602 723 605 746
rect 550 626 553 673
rect 546 623 553 626
rect 546 573 549 623
rect 554 576 557 616
rect 562 613 565 666
rect 562 583 565 606
rect 570 603 573 616
rect 578 593 581 606
rect 578 576 581 586
rect 554 573 581 576
rect 546 463 549 536
rect 554 533 557 573
rect 586 556 589 656
rect 594 603 597 616
rect 602 603 605 626
rect 610 603 613 646
rect 618 633 621 736
rect 618 593 621 606
rect 626 603 629 616
rect 634 603 637 763
rect 642 643 645 913
rect 650 903 653 1003
rect 658 1063 665 1066
rect 682 1103 693 1106
rect 658 976 661 1063
rect 682 1036 685 1103
rect 682 1033 693 1036
rect 698 1033 701 1086
rect 674 993 677 1016
rect 658 973 669 976
rect 666 933 669 973
rect 682 913 685 1006
rect 690 933 693 1033
rect 698 1003 701 1016
rect 650 723 653 806
rect 658 733 661 816
rect 666 793 669 816
rect 674 803 677 826
rect 682 803 685 816
rect 690 803 693 926
rect 650 603 653 636
rect 586 553 613 556
rect 554 513 557 526
rect 562 503 565 536
rect 554 473 573 476
rect 554 453 557 473
rect 562 446 565 466
rect 546 393 549 446
rect 554 443 565 446
rect 554 363 557 436
rect 570 426 573 473
rect 586 433 589 526
rect 562 413 565 426
rect 570 423 589 426
rect 570 413 581 416
rect 562 353 565 406
rect 570 403 581 406
rect 570 376 573 403
rect 570 373 581 376
rect 506 303 517 306
rect 530 293 533 326
rect 578 263 581 373
rect 586 363 589 423
rect 594 413 597 496
rect 610 443 613 553
rect 618 513 621 526
rect 626 523 629 556
rect 634 523 637 546
rect 642 533 645 586
rect 650 543 653 576
rect 666 556 669 766
rect 674 593 677 616
rect 682 586 685 796
rect 698 736 701 996
rect 706 966 709 1056
rect 722 1043 725 1126
rect 730 1106 733 1173
rect 738 1113 741 1146
rect 746 1133 749 1186
rect 754 1113 757 1196
rect 730 1103 749 1106
rect 706 963 713 966
rect 722 963 725 1006
rect 710 886 713 963
rect 738 936 741 1076
rect 746 1013 749 1103
rect 754 1016 757 1046
rect 770 1043 773 1336
rect 778 1276 781 1343
rect 786 1303 789 1326
rect 794 1306 797 1406
rect 802 1323 805 1416
rect 810 1373 813 1463
rect 818 1423 821 1456
rect 834 1436 837 1483
rect 826 1433 837 1436
rect 826 1403 829 1433
rect 834 1413 845 1416
rect 810 1316 813 1356
rect 826 1336 829 1366
rect 834 1343 837 1413
rect 842 1403 853 1406
rect 866 1403 869 1436
rect 818 1323 821 1336
rect 826 1333 845 1336
rect 850 1333 853 1396
rect 890 1393 893 1416
rect 914 1403 917 1573
rect 938 1566 941 1623
rect 946 1613 949 1734
rect 962 1693 965 1793
rect 970 1733 973 1746
rect 978 1733 981 1806
rect 986 1783 989 1813
rect 994 1733 997 1806
rect 1002 1743 1005 1816
rect 1010 1803 1013 1836
rect 1018 1736 1021 1876
rect 1026 1813 1029 1826
rect 1034 1813 1037 1856
rect 1010 1733 1021 1736
rect 994 1706 997 1726
rect 986 1703 997 1706
rect 986 1636 989 1703
rect 986 1633 997 1636
rect 954 1613 981 1616
rect 962 1583 965 1606
rect 930 1563 941 1566
rect 930 1533 933 1563
rect 930 1433 933 1526
rect 954 1513 957 1556
rect 978 1503 981 1526
rect 930 1423 957 1426
rect 866 1336 869 1386
rect 930 1366 933 1423
rect 922 1363 933 1366
rect 866 1333 873 1336
rect 810 1313 821 1316
rect 794 1303 801 1306
rect 778 1273 789 1276
rect 778 1183 781 1216
rect 786 1143 789 1273
rect 798 1236 801 1303
rect 794 1233 801 1236
rect 762 1023 773 1026
rect 754 1013 765 1016
rect 754 1003 765 1006
rect 770 953 773 1006
rect 778 1003 781 1136
rect 786 1003 789 1136
rect 794 1093 797 1233
rect 826 1226 829 1326
rect 842 1316 845 1333
rect 838 1313 845 1316
rect 850 1313 853 1326
rect 838 1236 841 1313
rect 838 1233 845 1236
rect 818 1223 829 1226
rect 802 1183 805 1216
rect 818 1203 821 1223
rect 826 1146 829 1216
rect 834 1193 837 1216
rect 842 1213 845 1233
rect 802 1123 805 1136
rect 810 1123 813 1146
rect 822 1143 829 1146
rect 802 1076 805 1116
rect 798 1073 805 1076
rect 798 1006 801 1073
rect 798 1003 805 1006
rect 786 983 789 996
rect 802 983 805 1003
rect 706 883 713 886
rect 706 866 709 883
rect 706 863 717 866
rect 706 853 709 863
rect 706 783 709 816
rect 714 813 717 863
rect 722 793 725 836
rect 730 776 733 936
rect 738 933 757 936
rect 658 553 669 556
rect 674 583 685 586
rect 690 733 701 736
rect 706 773 733 776
rect 674 553 677 583
rect 690 553 693 733
rect 698 703 701 726
rect 706 656 709 773
rect 714 733 717 766
rect 698 653 709 656
rect 698 556 701 653
rect 698 553 709 556
rect 642 463 645 526
rect 650 466 653 536
rect 658 533 661 553
rect 658 513 661 526
rect 650 463 661 466
rect 674 463 677 526
rect 602 413 605 426
rect 658 413 661 463
rect 682 413 685 516
rect 706 433 709 553
rect 714 533 717 726
rect 722 703 725 726
rect 730 723 733 766
rect 738 733 741 746
rect 738 713 741 726
rect 746 723 749 916
rect 754 896 757 926
rect 762 923 765 936
rect 778 933 781 946
rect 754 893 765 896
rect 762 836 765 893
rect 754 833 765 836
rect 754 773 757 833
rect 770 793 773 816
rect 754 733 757 746
rect 770 733 773 786
rect 778 776 781 926
rect 794 906 797 966
rect 810 933 813 1076
rect 822 1056 825 1143
rect 834 1123 837 1136
rect 834 1083 837 1116
rect 842 1076 845 1136
rect 850 1133 853 1306
rect 858 1213 861 1326
rect 870 1276 873 1333
rect 866 1273 873 1276
rect 866 1213 869 1273
rect 874 1213 877 1256
rect 850 1086 853 1126
rect 858 1093 861 1206
rect 882 1203 885 1216
rect 890 1196 893 1216
rect 898 1203 901 1276
rect 906 1213 909 1226
rect 914 1213 917 1326
rect 922 1286 925 1363
rect 938 1333 941 1376
rect 946 1353 949 1416
rect 954 1413 957 1423
rect 978 1413 981 1426
rect 954 1403 973 1406
rect 954 1333 957 1403
rect 986 1393 989 1616
rect 994 1613 997 1633
rect 994 1603 1005 1606
rect 1010 1583 1013 1733
rect 1018 1713 1021 1726
rect 1034 1723 1037 1766
rect 1026 1633 1029 1716
rect 994 1516 997 1536
rect 1018 1523 1021 1626
rect 1034 1613 1037 1646
rect 1042 1613 1045 1866
rect 1050 1623 1053 1896
rect 1066 1723 1069 1906
rect 1074 1733 1077 1816
rect 1074 1713 1077 1726
rect 1026 1603 1045 1606
rect 1050 1593 1053 1616
rect 1066 1605 1069 1646
rect 1034 1546 1037 1586
rect 1082 1556 1085 1886
rect 1178 1813 1181 1826
rect 1218 1813 1221 1836
rect 1226 1813 1229 1826
rect 1114 1766 1117 1806
rect 1138 1793 1141 1806
rect 1098 1763 1117 1766
rect 1090 1603 1093 1746
rect 1098 1593 1101 1763
rect 1114 1733 1117 1746
rect 1130 1733 1133 1756
rect 1154 1733 1157 1746
rect 1106 1613 1109 1626
rect 1114 1576 1117 1726
rect 1138 1703 1141 1726
rect 1194 1713 1197 1726
rect 1234 1723 1237 1816
rect 1242 1796 1245 1806
rect 1250 1803 1253 1856
rect 1258 1796 1261 1816
rect 1242 1793 1261 1796
rect 1242 1713 1245 1726
rect 1258 1683 1261 1726
rect 1146 1633 1165 1636
rect 1146 1613 1149 1633
rect 1154 1613 1157 1626
rect 1162 1603 1165 1633
rect 1170 1596 1173 1606
rect 1178 1603 1181 1656
rect 1266 1653 1269 1806
rect 1274 1793 1277 1940
rect 1298 1923 1301 1940
rect 1322 1906 1325 1926
rect 1314 1903 1325 1906
rect 1314 1836 1317 1903
rect 1314 1833 1325 1836
rect 1298 1803 1301 1816
rect 1274 1746 1277 1766
rect 1322 1763 1325 1833
rect 1330 1766 1333 1916
rect 1394 1913 1397 1940
rect 1338 1823 1341 1846
rect 1346 1813 1349 1836
rect 1330 1763 1341 1766
rect 1274 1743 1293 1746
rect 1290 1656 1293 1743
rect 1274 1653 1293 1656
rect 1186 1596 1189 1616
rect 1170 1593 1189 1596
rect 1114 1573 1125 1576
rect 1194 1573 1197 1606
rect 1066 1553 1085 1556
rect 1034 1543 1061 1546
rect 994 1513 1001 1516
rect 998 1436 1001 1513
rect 994 1433 1001 1436
rect 994 1413 997 1433
rect 1002 1403 1005 1416
rect 1010 1413 1013 1476
rect 1010 1356 1013 1406
rect 1026 1366 1029 1506
rect 1034 1453 1037 1543
rect 1042 1533 1053 1536
rect 1058 1533 1061 1543
rect 922 1283 933 1286
rect 906 1196 909 1206
rect 890 1193 909 1196
rect 914 1186 917 1206
rect 866 1133 869 1146
rect 882 1133 885 1186
rect 898 1183 917 1186
rect 866 1113 869 1126
rect 866 1086 869 1106
rect 850 1083 869 1086
rect 842 1073 853 1076
rect 818 1053 825 1056
rect 834 1056 837 1066
rect 834 1053 845 1056
rect 818 963 821 1053
rect 826 1013 829 1046
rect 834 1016 837 1026
rect 842 1023 845 1053
rect 834 1013 845 1016
rect 842 1003 845 1013
rect 850 1003 853 1073
rect 858 1003 861 1016
rect 818 923 821 946
rect 866 943 869 1016
rect 874 986 877 1026
rect 882 1013 885 1126
rect 898 1103 901 1183
rect 922 1166 925 1226
rect 930 1216 933 1283
rect 930 1213 941 1216
rect 914 1163 925 1166
rect 906 1123 909 1146
rect 882 996 885 1006
rect 890 1003 893 1026
rect 898 996 901 1016
rect 906 1003 909 1066
rect 914 1013 917 1163
rect 922 1023 925 1096
rect 882 993 901 996
rect 874 983 885 986
rect 914 983 917 1006
rect 846 933 869 936
rect 874 933 877 966
rect 882 933 885 983
rect 930 976 933 1206
rect 938 1173 941 1213
rect 946 1186 949 1216
rect 954 1213 957 1226
rect 962 1213 965 1356
rect 994 1353 1013 1356
rect 1018 1363 1029 1366
rect 970 1343 989 1346
rect 970 1323 973 1343
rect 978 1323 981 1336
rect 986 1333 989 1343
rect 994 1326 997 1353
rect 986 1323 997 1326
rect 986 1216 989 1323
rect 1002 1313 1005 1326
rect 962 1193 965 1206
rect 970 1196 973 1216
rect 978 1203 981 1216
rect 986 1213 997 1216
rect 1002 1213 1005 1226
rect 986 1196 989 1206
rect 970 1193 989 1196
rect 946 1183 965 1186
rect 914 973 933 976
rect 794 903 805 906
rect 802 846 805 903
rect 846 886 849 933
rect 858 916 861 926
rect 866 923 869 933
rect 874 916 877 926
rect 858 913 877 916
rect 890 906 893 926
rect 794 843 805 846
rect 842 883 849 886
rect 886 903 893 906
rect 778 773 789 776
rect 762 713 765 726
rect 754 663 765 666
rect 730 616 733 646
rect 722 613 733 616
rect 754 613 757 626
rect 762 616 765 663
rect 770 633 773 726
rect 786 723 789 773
rect 794 766 797 843
rect 810 783 813 806
rect 794 763 805 766
rect 762 613 773 616
rect 722 553 725 613
rect 730 603 741 606
rect 722 533 725 546
rect 730 533 733 603
rect 738 573 749 576
rect 714 443 717 526
rect 722 426 725 436
rect 706 423 725 426
rect 730 426 733 526
rect 738 493 741 573
rect 746 443 749 556
rect 754 533 757 586
rect 786 553 789 706
rect 802 603 805 763
rect 810 723 813 746
rect 818 576 821 816
rect 826 793 829 806
rect 834 803 837 816
rect 842 813 845 883
rect 886 836 889 903
rect 886 833 893 836
rect 858 803 861 816
rect 802 533 805 576
rect 810 573 821 576
rect 730 423 749 426
rect 706 413 709 423
rect 714 413 725 416
rect 594 393 597 406
rect 650 386 653 406
rect 658 393 661 406
rect 634 333 637 356
rect 474 233 477 256
rect 482 223 509 226
rect 514 223 525 226
rect 538 223 541 236
rect 554 233 581 236
rect 474 163 477 206
rect 482 183 485 223
rect 474 123 477 146
rect 410 96 413 106
rect 426 103 429 116
rect 410 93 429 96
rect 490 93 493 216
rect 498 193 501 206
rect 498 133 501 146
rect 506 143 509 186
rect 498 83 501 126
rect 506 123 509 136
rect 514 103 517 223
rect 522 213 549 216
rect 554 213 557 226
rect 562 213 565 226
rect 578 213 581 233
rect 586 213 589 326
rect 602 253 605 326
rect 618 286 621 326
rect 610 283 621 286
rect 610 213 613 283
rect 522 203 533 206
rect 522 163 525 203
rect 522 123 525 146
rect 578 133 581 176
rect 530 113 533 126
rect 546 93 549 126
rect 578 113 581 126
rect 586 83 589 186
rect 618 183 621 256
rect 634 253 637 326
rect 642 323 645 386
rect 650 383 661 386
rect 650 363 653 383
rect 666 253 669 326
rect 594 23 597 136
rect 602 123 605 136
rect 610 133 613 146
rect 626 133 629 206
rect 634 203 637 216
rect 642 203 645 216
rect 650 213 653 236
rect 666 213 669 226
rect 674 213 677 326
rect 690 296 693 386
rect 698 343 701 366
rect 706 326 709 396
rect 714 383 717 413
rect 722 356 725 406
rect 730 363 733 416
rect 738 383 741 416
rect 746 393 749 423
rect 754 413 757 526
rect 802 513 805 526
rect 810 506 813 573
rect 826 566 829 776
rect 842 766 845 796
rect 874 793 877 826
rect 890 813 893 833
rect 898 823 901 946
rect 906 933 909 946
rect 914 866 917 973
rect 938 966 941 1016
rect 946 1003 949 1026
rect 954 1013 957 1096
rect 962 1083 965 1183
rect 970 1133 973 1166
rect 994 1146 997 1213
rect 1018 1203 1021 1363
rect 1042 1336 1045 1526
rect 1050 1413 1053 1526
rect 1058 1423 1061 1526
rect 1066 1506 1069 1553
rect 1074 1543 1093 1546
rect 1074 1523 1077 1543
rect 1066 1503 1073 1506
rect 1070 1416 1073 1503
rect 1082 1473 1085 1536
rect 1090 1533 1093 1543
rect 1098 1486 1101 1536
rect 1106 1513 1109 1526
rect 1122 1503 1125 1573
rect 1146 1513 1149 1526
rect 1202 1523 1205 1536
rect 1210 1523 1213 1616
rect 1218 1543 1221 1626
rect 1250 1613 1253 1626
rect 1274 1606 1277 1653
rect 1282 1613 1285 1636
rect 1314 1633 1317 1716
rect 1274 1603 1285 1606
rect 1290 1603 1293 1616
rect 1314 1613 1317 1626
rect 1338 1603 1341 1763
rect 1346 1733 1349 1796
rect 1354 1753 1357 1816
rect 1362 1806 1365 1826
rect 1370 1813 1373 1836
rect 1362 1803 1373 1806
rect 1362 1733 1365 1746
rect 1386 1743 1389 1826
rect 1394 1813 1397 1906
rect 1394 1783 1397 1806
rect 1402 1803 1405 1816
rect 1410 1796 1413 1816
rect 1418 1803 1421 1856
rect 1426 1823 1429 1940
rect 1442 1903 1445 1940
rect 1506 1916 1509 1940
rect 1498 1913 1509 1916
rect 1498 1856 1501 1913
rect 1498 1853 1509 1856
rect 1426 1796 1429 1806
rect 1410 1793 1429 1796
rect 1434 1746 1437 1816
rect 1442 1813 1445 1826
rect 1482 1813 1485 1826
rect 1434 1743 1445 1746
rect 1346 1703 1349 1726
rect 1346 1603 1349 1696
rect 1386 1686 1389 1726
rect 1442 1723 1445 1743
rect 1450 1693 1453 1716
rect 1458 1713 1461 1806
rect 1290 1533 1293 1556
rect 1330 1533 1333 1546
rect 1338 1533 1341 1596
rect 1354 1556 1357 1686
rect 1370 1683 1389 1686
rect 1370 1613 1373 1683
rect 1378 1613 1381 1626
rect 1386 1603 1389 1656
rect 1394 1603 1397 1616
rect 1402 1573 1405 1606
rect 1410 1583 1413 1616
rect 1418 1613 1421 1626
rect 1346 1553 1357 1556
rect 1346 1526 1349 1553
rect 1378 1533 1381 1556
rect 1266 1513 1269 1526
rect 1306 1513 1309 1526
rect 1322 1523 1349 1526
rect 1362 1513 1365 1526
rect 1402 1513 1405 1526
rect 1458 1523 1461 1586
rect 1466 1533 1469 1606
rect 1474 1523 1477 1616
rect 1482 1503 1485 1806
rect 1506 1803 1509 1853
rect 1522 1816 1525 1906
rect 1690 1876 1693 1940
rect 1778 1937 1797 1940
rect 1690 1873 1701 1876
rect 1522 1813 1541 1816
rect 1522 1733 1525 1813
rect 1530 1733 1533 1806
rect 1554 1766 1557 1846
rect 1594 1803 1597 1816
rect 1554 1763 1581 1766
rect 1530 1716 1533 1726
rect 1538 1723 1541 1736
rect 1490 1703 1493 1716
rect 1498 1696 1501 1716
rect 1530 1713 1557 1716
rect 1578 1706 1581 1763
rect 1602 1713 1605 1726
rect 1570 1703 1581 1706
rect 1498 1693 1509 1696
rect 1506 1646 1509 1693
rect 1498 1643 1509 1646
rect 1498 1593 1501 1643
rect 1562 1613 1565 1626
rect 1522 1583 1525 1606
rect 1562 1533 1565 1596
rect 1570 1583 1573 1703
rect 1610 1623 1613 1726
rect 1626 1656 1629 1726
rect 1634 1723 1637 1736
rect 1642 1723 1645 1806
rect 1626 1653 1637 1656
rect 1602 1553 1605 1616
rect 1618 1613 1629 1616
rect 1634 1613 1637 1653
rect 1650 1626 1653 1856
rect 1658 1796 1661 1816
rect 1666 1803 1669 1816
rect 1682 1806 1685 1816
rect 1690 1813 1693 1826
rect 1698 1806 1701 1873
rect 1738 1813 1741 1826
rect 1674 1796 1677 1806
rect 1682 1803 1701 1806
rect 1658 1793 1677 1796
rect 1746 1736 1749 1806
rect 1658 1683 1661 1726
rect 1714 1713 1717 1736
rect 1738 1733 1749 1736
rect 1754 1733 1757 1756
rect 1738 1713 1741 1733
rect 1746 1673 1749 1726
rect 1762 1696 1765 1816
rect 1778 1773 1781 1806
rect 1794 1736 1797 1937
rect 1802 1803 1805 1816
rect 1810 1796 1813 1816
rect 1818 1803 1821 1856
rect 1834 1813 1837 1826
rect 1826 1796 1829 1806
rect 1810 1793 1829 1796
rect 1758 1693 1765 1696
rect 1778 1696 1781 1736
rect 1786 1733 1797 1736
rect 1786 1713 1789 1733
rect 1778 1693 1789 1696
rect 1758 1646 1761 1693
rect 1758 1643 1765 1646
rect 1642 1623 1653 1626
rect 1618 1593 1621 1606
rect 1626 1603 1629 1613
rect 1594 1543 1613 1546
rect 1594 1533 1597 1543
rect 1538 1513 1541 1526
rect 1578 1513 1581 1526
rect 1586 1503 1589 1526
rect 1602 1523 1605 1536
rect 1610 1523 1613 1543
rect 1618 1533 1621 1576
rect 1642 1573 1645 1623
rect 1650 1566 1653 1616
rect 1706 1613 1709 1626
rect 1666 1583 1669 1606
rect 1650 1563 1669 1566
rect 1626 1523 1629 1556
rect 1642 1533 1645 1546
rect 1666 1523 1669 1563
rect 1730 1533 1733 1576
rect 1746 1533 1749 1616
rect 1754 1613 1757 1626
rect 1762 1606 1765 1643
rect 1770 1613 1773 1686
rect 1786 1616 1789 1693
rect 1778 1613 1789 1616
rect 1754 1603 1765 1606
rect 1746 1506 1749 1526
rect 1754 1513 1757 1603
rect 1738 1503 1749 1506
rect 1098 1483 1109 1486
rect 1106 1426 1109 1483
rect 1738 1446 1741 1503
rect 1106 1423 1125 1426
rect 1066 1413 1073 1416
rect 1098 1413 1109 1416
rect 1050 1386 1053 1406
rect 1050 1383 1057 1386
rect 1034 1333 1045 1336
rect 1034 1193 1037 1333
rect 1042 1313 1045 1325
rect 1054 1306 1057 1383
rect 1066 1353 1069 1413
rect 1050 1303 1057 1306
rect 1042 1213 1045 1226
rect 978 1143 997 1146
rect 978 1123 981 1143
rect 986 1133 997 1136
rect 970 1016 973 1116
rect 986 1056 989 1133
rect 978 1053 989 1056
rect 978 1023 981 1053
rect 954 983 957 1006
rect 922 963 941 966
rect 922 923 925 963
rect 930 873 933 946
rect 938 923 941 936
rect 938 886 941 916
rect 946 893 949 956
rect 954 923 957 966
rect 962 933 965 1016
rect 970 1013 981 1016
rect 986 1013 989 1026
rect 994 1013 997 1126
rect 1002 1023 1005 1046
rect 1010 1016 1013 1176
rect 1050 1173 1053 1303
rect 1082 1206 1085 1366
rect 1106 1333 1109 1413
rect 1114 1363 1117 1416
rect 1122 1413 1125 1423
rect 1130 1346 1133 1406
rect 1114 1343 1133 1346
rect 1090 1323 1101 1326
rect 1098 1266 1101 1323
rect 1106 1273 1109 1326
rect 1114 1316 1117 1343
rect 1130 1323 1133 1336
rect 1138 1326 1141 1416
rect 1146 1333 1149 1366
rect 1154 1343 1157 1426
rect 1194 1413 1197 1436
rect 1234 1413 1253 1416
rect 1274 1413 1277 1426
rect 1298 1413 1301 1426
rect 1322 1413 1341 1416
rect 1346 1413 1349 1436
rect 1362 1413 1365 1426
rect 1378 1413 1381 1436
rect 1386 1413 1397 1416
rect 1402 1413 1405 1426
rect 1426 1413 1445 1416
rect 1466 1413 1469 1436
rect 1530 1413 1533 1426
rect 1562 1413 1565 1446
rect 1738 1443 1749 1446
rect 1170 1333 1173 1346
rect 1138 1323 1149 1326
rect 1114 1313 1125 1316
rect 1098 1263 1109 1266
rect 1098 1216 1101 1236
rect 1090 1213 1101 1216
rect 1106 1213 1109 1263
rect 1122 1253 1125 1313
rect 1082 1203 1101 1206
rect 1098 1133 1101 1203
rect 1114 1173 1117 1216
rect 1122 1213 1125 1236
rect 1130 1196 1133 1276
rect 1138 1213 1141 1236
rect 1146 1213 1149 1256
rect 1162 1226 1165 1236
rect 1154 1223 1165 1226
rect 1154 1213 1157 1223
rect 1138 1203 1149 1206
rect 1130 1193 1141 1196
rect 1050 1123 1061 1126
rect 1098 1083 1101 1126
rect 1106 1123 1109 1156
rect 1114 1123 1117 1136
rect 1002 1013 1013 1016
rect 1018 1053 1037 1056
rect 954 903 957 916
rect 938 883 949 886
rect 914 863 925 866
rect 802 503 813 506
rect 818 563 829 566
rect 834 763 845 766
rect 770 413 773 426
rect 786 413 789 466
rect 802 413 805 503
rect 818 496 821 563
rect 826 503 829 526
rect 810 493 821 496
rect 810 413 813 493
rect 754 356 757 406
rect 818 376 821 406
rect 722 353 757 356
rect 714 333 717 346
rect 770 333 773 346
rect 706 323 717 326
rect 686 293 693 296
rect 686 226 689 293
rect 686 223 693 226
rect 658 203 677 206
rect 690 203 693 223
rect 674 193 677 203
rect 698 196 701 316
rect 722 276 725 326
rect 778 313 781 376
rect 786 373 821 376
rect 786 333 789 373
rect 786 303 789 326
rect 794 323 797 366
rect 826 356 829 416
rect 802 353 829 356
rect 802 276 805 353
rect 810 343 829 346
rect 834 343 837 763
rect 842 613 845 626
rect 842 523 845 606
rect 866 576 869 746
rect 874 733 877 756
rect 874 613 877 646
rect 882 633 885 806
rect 898 793 901 816
rect 890 623 893 736
rect 898 643 901 726
rect 906 696 909 786
rect 914 733 917 746
rect 914 713 917 726
rect 906 693 913 696
rect 850 573 869 576
rect 882 573 885 616
rect 898 613 901 636
rect 910 626 913 693
rect 922 683 925 863
rect 930 633 933 846
rect 938 813 941 856
rect 946 823 949 883
rect 962 826 965 926
rect 970 916 973 1006
rect 978 1003 981 1013
rect 986 996 989 1006
rect 978 993 989 996
rect 978 923 981 993
rect 970 913 981 916
rect 986 833 989 986
rect 1002 963 1005 1013
rect 1010 983 1013 1006
rect 1018 953 1021 1053
rect 1034 1046 1037 1053
rect 1026 1023 1029 1046
rect 1034 1043 1045 1046
rect 1050 1043 1069 1046
rect 1050 1036 1053 1043
rect 1042 1033 1053 1036
rect 1042 1023 1053 1026
rect 1026 1013 1037 1016
rect 1034 956 1037 1013
rect 1050 983 1053 1016
rect 1058 1013 1061 1036
rect 1066 963 1069 1043
rect 1074 1003 1077 1026
rect 1098 1013 1101 1046
rect 1106 1013 1109 1106
rect 1122 1003 1125 1126
rect 1130 1113 1133 1146
rect 1138 1133 1141 1193
rect 1146 1113 1149 1156
rect 1162 1153 1165 1216
rect 1178 1213 1181 1226
rect 1186 1213 1189 1366
rect 1194 1323 1197 1336
rect 1202 1273 1205 1356
rect 1242 1353 1245 1406
rect 1250 1363 1253 1413
rect 1298 1393 1301 1406
rect 1306 1373 1309 1406
rect 1330 1393 1333 1406
rect 1266 1333 1269 1346
rect 1314 1333 1333 1336
rect 1210 1266 1213 1326
rect 1234 1323 1245 1326
rect 1202 1263 1213 1266
rect 1170 1193 1173 1206
rect 1154 1133 1165 1136
rect 1170 1133 1173 1146
rect 1178 1133 1181 1176
rect 1186 1143 1189 1206
rect 1194 1153 1197 1206
rect 1202 1203 1205 1263
rect 1258 1253 1261 1326
rect 1314 1303 1317 1326
rect 1218 1176 1221 1206
rect 1130 1003 1133 1016
rect 1138 1013 1141 1026
rect 1138 996 1141 1006
rect 1146 1003 1149 1046
rect 1154 1033 1157 1066
rect 1162 1056 1165 1126
rect 1178 1113 1181 1126
rect 1186 1106 1189 1126
rect 1194 1113 1197 1136
rect 1202 1123 1205 1176
rect 1218 1173 1229 1176
rect 1210 1133 1213 1146
rect 1226 1133 1229 1173
rect 1234 1166 1237 1216
rect 1242 1193 1245 1216
rect 1282 1166 1285 1216
rect 1234 1163 1245 1166
rect 1178 1103 1189 1106
rect 1178 1056 1181 1066
rect 1162 1053 1181 1056
rect 1162 1023 1173 1026
rect 1154 1013 1173 1016
rect 1154 1003 1173 1006
rect 1178 1003 1181 1053
rect 1186 1003 1189 1016
rect 1154 996 1157 1003
rect 1138 993 1157 996
rect 1034 953 1045 956
rect 1010 883 1013 926
rect 962 823 989 826
rect 946 803 949 816
rect 954 803 957 816
rect 962 793 965 806
rect 970 756 973 816
rect 986 813 989 823
rect 1002 813 1005 866
rect 1034 813 1037 926
rect 1042 903 1045 953
rect 1050 933 1053 956
rect 1042 823 1045 836
rect 1050 808 1053 926
rect 1058 813 1061 926
rect 1082 923 1093 926
rect 1066 813 1069 866
rect 978 783 981 806
rect 986 766 989 806
rect 1034 805 1053 808
rect 986 763 1005 766
rect 970 753 981 756
rect 946 713 949 726
rect 978 723 981 753
rect 986 733 989 746
rect 910 623 925 626
rect 850 503 853 573
rect 890 563 893 606
rect 906 593 909 606
rect 914 556 917 616
rect 922 603 925 623
rect 938 603 941 666
rect 954 583 957 686
rect 962 593 965 616
rect 898 553 917 556
rect 898 533 901 553
rect 906 533 909 546
rect 882 513 885 526
rect 898 513 901 526
rect 842 433 877 436
rect 810 323 813 343
rect 818 323 821 336
rect 826 333 829 343
rect 842 336 845 433
rect 850 413 853 426
rect 874 413 877 433
rect 882 413 885 426
rect 850 376 853 406
rect 850 373 861 376
rect 834 333 845 336
rect 826 313 829 326
rect 706 273 725 276
rect 794 273 805 276
rect 706 213 709 273
rect 682 193 701 196
rect 674 133 677 186
rect 618 103 621 126
rect 626 113 629 126
rect 682 73 685 193
rect 722 183 725 236
rect 730 213 733 226
rect 738 223 757 226
rect 762 223 773 226
rect 738 213 749 216
rect 730 133 733 206
rect 746 193 749 206
rect 738 126 741 166
rect 730 123 741 126
rect 746 123 749 186
rect 754 173 757 223
rect 778 213 781 266
rect 786 213 789 246
rect 762 13 765 136
rect 770 133 773 206
rect 778 203 789 206
rect 794 193 797 273
rect 802 173 805 216
rect 810 156 813 206
rect 818 203 821 306
rect 826 233 829 296
rect 826 203 829 216
rect 834 183 837 333
rect 842 283 845 326
rect 858 283 861 346
rect 898 336 901 416
rect 906 403 909 526
rect 914 433 917 496
rect 938 413 941 526
rect 954 413 957 546
rect 962 523 965 556
rect 970 543 973 646
rect 986 643 989 726
rect 994 713 997 756
rect 1002 723 1005 763
rect 1010 696 1013 736
rect 1018 733 1021 766
rect 1010 693 1021 696
rect 978 563 981 626
rect 986 573 989 596
rect 1002 573 1005 636
rect 1010 556 1013 686
rect 1018 603 1021 693
rect 1026 663 1029 786
rect 1058 763 1061 806
rect 1074 803 1085 806
rect 1074 733 1077 796
rect 1090 786 1093 826
rect 1106 823 1109 866
rect 1098 805 1101 816
rect 1114 796 1117 946
rect 1122 903 1125 986
rect 1194 946 1197 1106
rect 1242 1103 1245 1163
rect 1274 1163 1285 1166
rect 1266 1136 1269 1156
rect 1262 1133 1269 1136
rect 1250 1113 1253 1126
rect 1262 1056 1265 1133
rect 1210 1036 1213 1056
rect 1242 1036 1245 1056
rect 1262 1053 1269 1056
rect 1210 1033 1245 1036
rect 1202 1013 1205 1026
rect 1210 1013 1213 1033
rect 1218 1006 1221 1026
rect 1234 1013 1237 1026
rect 1202 983 1205 1006
rect 1210 1003 1221 1006
rect 1226 1003 1237 1006
rect 1242 1003 1245 1033
rect 1258 1026 1261 1036
rect 1250 1023 1261 1026
rect 1250 1003 1261 1006
rect 1258 976 1261 996
rect 1266 983 1269 1053
rect 1274 1036 1277 1163
rect 1290 1153 1293 1286
rect 1322 1283 1325 1326
rect 1330 1276 1333 1333
rect 1338 1323 1341 1413
rect 1346 1343 1349 1406
rect 1354 1373 1357 1406
rect 1346 1326 1349 1336
rect 1354 1333 1357 1356
rect 1346 1323 1357 1326
rect 1362 1303 1365 1336
rect 1370 1333 1373 1406
rect 1314 1273 1333 1276
rect 1298 1183 1301 1216
rect 1306 1193 1309 1206
rect 1314 1203 1317 1273
rect 1322 1186 1325 1256
rect 1330 1213 1333 1226
rect 1346 1213 1349 1276
rect 1370 1253 1373 1326
rect 1378 1213 1381 1386
rect 1386 1333 1389 1406
rect 1394 1383 1397 1413
rect 1410 1393 1413 1406
rect 1418 1376 1421 1406
rect 1394 1373 1421 1376
rect 1386 1293 1389 1326
rect 1394 1266 1397 1373
rect 1410 1313 1413 1326
rect 1442 1306 1445 1413
rect 1498 1376 1501 1406
rect 1474 1373 1501 1376
rect 1450 1333 1453 1346
rect 1474 1333 1477 1373
rect 1482 1336 1485 1346
rect 1482 1333 1493 1336
rect 1506 1333 1509 1406
rect 1514 1333 1517 1346
rect 1458 1323 1477 1326
rect 1434 1303 1445 1306
rect 1394 1263 1413 1266
rect 1330 1193 1333 1206
rect 1322 1183 1333 1186
rect 1314 1133 1317 1146
rect 1306 1113 1309 1126
rect 1274 1033 1285 1036
rect 1282 1023 1285 1033
rect 1298 1013 1301 1066
rect 1314 1013 1317 1126
rect 1314 993 1317 1006
rect 1258 973 1269 976
rect 1146 943 1165 946
rect 1130 876 1133 926
rect 1138 886 1141 936
rect 1146 933 1149 943
rect 1146 893 1149 926
rect 1138 883 1149 886
rect 1130 873 1141 876
rect 1122 823 1125 836
rect 1138 823 1141 873
rect 1146 823 1149 883
rect 1122 813 1149 816
rect 1122 803 1133 806
rect 1114 793 1133 796
rect 1090 783 1125 786
rect 1122 773 1125 783
rect 1050 693 1053 726
rect 1026 613 1029 646
rect 1058 623 1061 716
rect 1074 693 1077 726
rect 1066 653 1069 686
rect 1026 596 1029 606
rect 1074 603 1077 666
rect 1082 653 1085 726
rect 1106 723 1117 726
rect 1130 713 1133 793
rect 1138 663 1141 766
rect 1146 743 1149 776
rect 1154 733 1157 936
rect 1162 933 1165 943
rect 1178 943 1197 946
rect 1162 893 1165 926
rect 1170 923 1173 936
rect 1162 753 1165 836
rect 1178 833 1181 943
rect 1186 903 1189 926
rect 1194 813 1197 936
rect 1210 933 1213 946
rect 1202 923 1213 926
rect 1218 923 1221 936
rect 1226 883 1229 926
rect 1234 903 1237 936
rect 1242 933 1253 936
rect 1258 933 1261 966
rect 1266 956 1269 973
rect 1282 963 1285 986
rect 1290 983 1301 986
rect 1290 956 1293 983
rect 1322 976 1325 1156
rect 1330 1123 1333 1183
rect 1338 1133 1341 1186
rect 1346 1086 1349 1146
rect 1362 1133 1365 1166
rect 1378 1143 1381 1206
rect 1386 1136 1389 1216
rect 1402 1213 1405 1256
rect 1386 1133 1397 1136
rect 1378 1123 1389 1126
rect 1394 1116 1397 1133
rect 1394 1113 1401 1116
rect 1346 1083 1357 1086
rect 1354 1013 1357 1083
rect 1378 1013 1381 1046
rect 1266 953 1293 956
rect 1314 973 1325 976
rect 1266 936 1269 946
rect 1298 943 1309 946
rect 1266 933 1277 936
rect 1242 863 1245 926
rect 1266 906 1269 926
rect 1258 903 1269 906
rect 1258 846 1261 903
rect 1258 843 1269 846
rect 1274 843 1277 933
rect 1282 903 1285 926
rect 1298 923 1301 943
rect 1314 936 1317 973
rect 1306 933 1317 936
rect 1290 873 1293 916
rect 1306 903 1309 933
rect 1314 883 1317 916
rect 1322 903 1325 916
rect 1330 903 1333 966
rect 1338 893 1341 926
rect 1346 923 1349 946
rect 1346 903 1349 916
rect 1354 913 1357 956
rect 1362 903 1365 986
rect 1370 936 1373 1006
rect 1378 983 1381 1006
rect 1370 933 1381 936
rect 1386 933 1389 1086
rect 1398 1046 1401 1113
rect 1410 1103 1413 1263
rect 1426 1203 1429 1226
rect 1434 1146 1437 1303
rect 1474 1256 1477 1316
rect 1466 1253 1477 1256
rect 1458 1223 1461 1236
rect 1466 1216 1469 1253
rect 1482 1223 1485 1326
rect 1490 1316 1493 1333
rect 1490 1313 1497 1316
rect 1494 1226 1497 1313
rect 1506 1233 1509 1316
rect 1514 1263 1517 1325
rect 1522 1273 1525 1336
rect 1530 1333 1541 1336
rect 1546 1333 1549 1346
rect 1554 1333 1557 1406
rect 1562 1333 1565 1406
rect 1578 1393 1581 1416
rect 1490 1223 1497 1226
rect 1530 1223 1533 1326
rect 1538 1323 1549 1326
rect 1538 1243 1541 1323
rect 1554 1322 1565 1325
rect 1570 1323 1573 1356
rect 1546 1313 1557 1316
rect 1546 1296 1549 1313
rect 1546 1293 1553 1296
rect 1562 1293 1565 1322
rect 1550 1226 1553 1293
rect 1578 1283 1581 1366
rect 1586 1333 1589 1416
rect 1602 1413 1605 1426
rect 1634 1413 1637 1426
rect 1674 1413 1693 1416
rect 1714 1413 1717 1426
rect 1594 1363 1597 1406
rect 1602 1383 1605 1406
rect 1594 1333 1613 1336
rect 1594 1313 1597 1326
rect 1546 1223 1553 1226
rect 1442 1213 1469 1216
rect 1490 1206 1493 1223
rect 1466 1203 1493 1206
rect 1430 1143 1437 1146
rect 1430 1086 1433 1143
rect 1442 1093 1445 1196
rect 1466 1153 1469 1203
rect 1506 1193 1517 1196
rect 1506 1163 1509 1186
rect 1450 1133 1453 1146
rect 1474 1103 1477 1126
rect 1498 1096 1501 1156
rect 1506 1133 1509 1146
rect 1506 1103 1509 1126
rect 1514 1116 1517 1136
rect 1522 1123 1525 1206
rect 1530 1203 1533 1216
rect 1538 1143 1541 1216
rect 1546 1193 1549 1223
rect 1586 1213 1589 1306
rect 1602 1233 1605 1333
rect 1610 1323 1621 1326
rect 1610 1213 1613 1323
rect 1634 1316 1637 1336
rect 1642 1333 1645 1386
rect 1674 1356 1677 1413
rect 1658 1353 1677 1356
rect 1682 1396 1685 1406
rect 1682 1393 1693 1396
rect 1738 1393 1741 1406
rect 1746 1403 1749 1443
rect 1762 1433 1765 1596
rect 1778 1593 1781 1613
rect 1770 1533 1773 1576
rect 1770 1513 1773 1526
rect 1778 1456 1781 1566
rect 1786 1523 1789 1536
rect 1794 1533 1797 1576
rect 1802 1563 1805 1776
rect 1842 1723 1845 1816
rect 1858 1793 1861 1806
rect 1866 1733 1869 1776
rect 1882 1723 1885 1816
rect 1938 1813 1941 1826
rect 1834 1623 1861 1626
rect 1850 1603 1853 1616
rect 1858 1613 1861 1623
rect 1802 1543 1821 1546
rect 1802 1523 1805 1543
rect 1810 1513 1813 1536
rect 1818 1533 1821 1543
rect 1826 1523 1829 1596
rect 1858 1593 1861 1606
rect 1866 1603 1869 1716
rect 1898 1683 1901 1726
rect 1890 1623 1893 1676
rect 1930 1623 1933 1736
rect 1858 1533 1861 1566
rect 1842 1513 1845 1526
rect 1882 1513 1885 1526
rect 1938 1523 1941 1596
rect 1770 1453 1781 1456
rect 1754 1413 1757 1426
rect 1770 1403 1773 1453
rect 1794 1413 1797 1426
rect 1850 1413 1853 1506
rect 1658 1326 1661 1353
rect 1666 1333 1669 1346
rect 1682 1336 1685 1393
rect 1674 1333 1685 1336
rect 1738 1333 1741 1346
rect 1858 1336 1861 1406
rect 1658 1323 1669 1326
rect 1626 1313 1645 1316
rect 1650 1276 1653 1316
rect 1642 1273 1653 1276
rect 1554 1153 1557 1206
rect 1562 1193 1565 1206
rect 1610 1183 1613 1206
rect 1514 1113 1525 1116
rect 1530 1113 1533 1136
rect 1490 1093 1501 1096
rect 1394 1043 1401 1046
rect 1426 1083 1433 1086
rect 1394 1013 1397 1043
rect 1426 1013 1429 1083
rect 1442 1013 1445 1066
rect 1490 1036 1493 1093
rect 1506 1073 1517 1076
rect 1522 1073 1525 1113
rect 1450 1033 1469 1036
rect 1394 963 1397 1006
rect 1378 926 1381 933
rect 1370 863 1373 926
rect 1378 923 1389 926
rect 1378 903 1381 916
rect 1386 906 1389 923
rect 1386 903 1405 906
rect 1162 733 1165 746
rect 1170 733 1173 766
rect 1210 763 1213 836
rect 1218 813 1221 826
rect 1242 813 1245 826
rect 1218 773 1221 806
rect 1266 753 1269 843
rect 1274 813 1277 826
rect 1274 773 1277 806
rect 1282 783 1285 836
rect 1290 803 1293 816
rect 1298 773 1301 856
rect 1306 813 1309 846
rect 1314 813 1317 826
rect 1330 813 1333 846
rect 1362 813 1365 846
rect 1394 813 1397 826
rect 1402 813 1405 903
rect 1418 846 1421 926
rect 1418 843 1429 846
rect 1418 813 1421 826
rect 1306 783 1309 806
rect 1314 773 1317 806
rect 1154 723 1173 726
rect 1098 613 1101 626
rect 1082 596 1085 606
rect 1130 603 1133 636
rect 978 553 1013 556
rect 1018 593 1029 596
rect 1074 593 1085 596
rect 1018 553 1021 593
rect 978 533 981 553
rect 1026 533 1029 566
rect 1074 553 1077 593
rect 970 516 973 526
rect 962 513 973 516
rect 970 493 973 513
rect 954 383 957 406
rect 890 333 901 336
rect 842 213 845 256
rect 850 213 853 226
rect 866 213 869 226
rect 850 193 853 206
rect 810 153 821 156
rect 818 133 821 153
rect 826 133 829 166
rect 858 163 861 206
rect 874 203 877 306
rect 882 203 885 316
rect 890 293 893 333
rect 890 223 893 276
rect 898 263 901 326
rect 906 313 909 326
rect 906 233 909 276
rect 874 133 877 186
rect 890 183 893 216
rect 898 213 901 226
rect 914 223 917 286
rect 922 203 925 316
rect 930 303 933 326
rect 938 313 941 326
rect 954 316 957 336
rect 962 333 965 426
rect 978 413 981 526
rect 986 406 989 506
rect 994 413 997 426
rect 1010 413 1013 526
rect 1026 513 1029 526
rect 1034 503 1037 536
rect 1090 533 1093 556
rect 1106 533 1117 536
rect 1026 466 1029 476
rect 1026 463 1061 466
rect 1018 413 1021 426
rect 970 393 973 406
rect 978 353 981 406
rect 986 403 997 406
rect 994 373 997 403
rect 1002 353 1005 406
rect 1010 333 1013 406
rect 1026 353 1029 436
rect 1042 413 1053 416
rect 1074 413 1077 506
rect 1082 413 1085 526
rect 1098 503 1101 526
rect 1106 513 1109 526
rect 1034 363 1037 406
rect 1042 396 1045 413
rect 1050 403 1061 406
rect 1042 393 1053 396
rect 1050 376 1053 393
rect 1058 386 1061 403
rect 1066 393 1069 406
rect 1058 383 1069 386
rect 1074 383 1077 406
rect 1050 373 1061 376
rect 1066 333 1069 383
rect 1074 333 1077 376
rect 1090 353 1093 456
rect 1106 436 1109 456
rect 1098 433 1109 436
rect 1098 413 1101 426
rect 1114 413 1117 526
rect 1098 393 1101 406
rect 1106 403 1117 406
rect 1106 373 1109 403
rect 1122 363 1125 576
rect 1130 533 1133 586
rect 1138 533 1141 626
rect 1154 613 1157 723
rect 1194 713 1197 726
rect 1186 613 1189 656
rect 1122 333 1125 346
rect 954 313 961 316
rect 930 213 933 226
rect 882 143 885 166
rect 938 133 941 296
rect 946 196 949 306
rect 958 246 961 313
rect 978 303 981 326
rect 954 243 961 246
rect 954 223 957 243
rect 970 213 973 256
rect 1018 246 1021 326
rect 1042 313 1045 326
rect 1018 243 1045 246
rect 1002 233 1013 236
rect 1002 223 1005 233
rect 1010 213 1013 226
rect 1018 213 1021 226
rect 946 193 957 196
rect 1002 193 1005 206
rect 954 156 957 193
rect 954 153 965 156
rect 946 133 949 146
rect 770 113 773 126
rect 794 123 805 126
rect 818 113 821 126
rect 850 113 853 126
rect 882 93 885 126
rect 906 103 909 126
rect 954 83 957 126
rect 962 43 965 153
rect 970 63 973 186
rect 986 156 989 186
rect 978 153 989 156
rect 978 143 981 153
rect 978 113 981 126
rect 1026 123 1029 236
rect 1042 213 1045 243
rect 1050 213 1053 326
rect 1106 236 1109 326
rect 1130 323 1133 516
rect 1138 493 1141 516
rect 1146 473 1149 586
rect 1186 583 1189 606
rect 1170 546 1173 566
rect 1154 543 1173 546
rect 1154 523 1157 543
rect 1162 493 1165 536
rect 1170 533 1173 543
rect 1170 503 1173 526
rect 1178 506 1181 536
rect 1186 516 1189 556
rect 1194 523 1197 626
rect 1202 583 1205 666
rect 1218 633 1221 746
rect 1298 743 1325 746
rect 1234 733 1245 736
rect 1210 553 1213 616
rect 1226 613 1229 726
rect 1234 686 1237 726
rect 1242 706 1245 726
rect 1274 713 1277 726
rect 1290 723 1293 736
rect 1306 713 1309 736
rect 1314 723 1317 736
rect 1322 733 1325 743
rect 1330 713 1333 746
rect 1346 733 1349 766
rect 1362 743 1365 796
rect 1370 736 1373 806
rect 1362 733 1381 736
rect 1386 733 1389 786
rect 1418 783 1421 806
rect 1338 723 1349 726
rect 1242 703 1253 706
rect 1234 683 1241 686
rect 1238 606 1241 683
rect 1218 563 1221 606
rect 1234 603 1241 606
rect 1250 603 1253 703
rect 1234 553 1237 603
rect 1186 513 1197 516
rect 1178 503 1189 506
rect 1138 436 1141 466
rect 1154 443 1157 466
rect 1186 456 1189 503
rect 1178 453 1189 456
rect 1138 433 1157 436
rect 1138 413 1141 426
rect 1154 423 1157 433
rect 1170 413 1173 446
rect 1186 413 1189 453
rect 1194 413 1197 456
rect 1138 303 1141 356
rect 1146 353 1157 356
rect 1146 296 1149 353
rect 1130 293 1149 296
rect 1090 233 1109 236
rect 1058 223 1077 226
rect 1090 216 1093 233
rect 1074 213 1093 216
rect 1098 213 1101 226
rect 1106 223 1109 233
rect 1122 223 1125 236
rect 1050 203 1069 206
rect 1034 133 1037 146
rect 1034 93 1037 126
rect 1042 73 1045 136
rect 1050 123 1053 203
rect 1074 193 1077 206
rect 1090 203 1125 206
rect 1058 33 1061 136
rect 1066 123 1069 146
rect 1074 133 1077 166
rect 1122 133 1125 196
rect 1082 0 1085 16
rect 1098 0 1101 76
rect 1122 73 1125 126
rect 1130 13 1133 293
rect 1138 233 1141 266
rect 1154 223 1157 346
rect 1162 223 1165 376
rect 1178 356 1181 376
rect 1174 353 1181 356
rect 1186 353 1189 406
rect 1174 236 1177 353
rect 1194 336 1197 406
rect 1202 373 1205 546
rect 1250 533 1253 546
rect 1258 533 1261 706
rect 1266 633 1269 646
rect 1274 623 1277 636
rect 1266 603 1277 606
rect 1282 586 1285 626
rect 1290 603 1293 616
rect 1314 613 1317 636
rect 1322 613 1325 696
rect 1346 656 1349 723
rect 1354 673 1357 726
rect 1362 706 1365 733
rect 1370 713 1373 726
rect 1362 703 1373 706
rect 1346 653 1365 656
rect 1282 583 1309 586
rect 1218 506 1221 526
rect 1210 503 1221 506
rect 1210 443 1213 503
rect 1210 343 1213 416
rect 1218 403 1221 486
rect 1234 456 1237 516
rect 1258 513 1261 526
rect 1282 503 1285 526
rect 1290 513 1293 526
rect 1306 483 1309 583
rect 1314 516 1317 586
rect 1322 533 1325 556
rect 1330 523 1333 536
rect 1314 513 1333 516
rect 1234 453 1301 456
rect 1226 403 1229 446
rect 1250 443 1285 446
rect 1250 436 1253 443
rect 1234 433 1253 436
rect 1234 413 1237 433
rect 1250 423 1261 426
rect 1258 413 1261 423
rect 1266 413 1269 426
rect 1282 423 1285 443
rect 1298 413 1301 453
rect 1306 413 1309 446
rect 1314 406 1317 506
rect 1322 433 1325 486
rect 1330 416 1333 513
rect 1234 396 1237 406
rect 1282 403 1317 406
rect 1322 413 1333 416
rect 1338 416 1341 646
rect 1346 533 1349 626
rect 1354 593 1357 616
rect 1362 613 1365 653
rect 1362 553 1365 606
rect 1370 563 1373 703
rect 1378 613 1381 726
rect 1378 596 1381 606
rect 1386 603 1389 676
rect 1394 613 1397 766
rect 1426 753 1429 843
rect 1434 833 1437 936
rect 1442 933 1445 1006
rect 1450 943 1453 1033
rect 1466 1013 1469 1033
rect 1482 1033 1493 1036
rect 1482 1013 1485 1033
rect 1498 1013 1501 1026
rect 1506 1013 1509 1066
rect 1498 986 1501 1006
rect 1490 983 1501 986
rect 1458 936 1461 966
rect 1450 933 1461 936
rect 1466 933 1469 956
rect 1490 943 1493 983
rect 1506 973 1509 1006
rect 1514 976 1517 1073
rect 1530 1066 1533 1086
rect 1538 1076 1541 1126
rect 1546 1103 1549 1126
rect 1538 1073 1549 1076
rect 1530 1063 1541 1066
rect 1522 1003 1525 1056
rect 1538 1053 1541 1063
rect 1546 1013 1549 1073
rect 1554 1023 1557 1086
rect 1570 1006 1573 1016
rect 1578 1013 1581 1026
rect 1586 1013 1589 1056
rect 1594 1013 1597 1156
rect 1602 1133 1605 1176
rect 1602 1006 1605 1126
rect 1610 1066 1613 1136
rect 1618 1123 1621 1236
rect 1642 1223 1645 1273
rect 1666 1213 1669 1323
rect 1674 1223 1677 1333
rect 1682 1306 1685 1326
rect 1706 1323 1717 1326
rect 1730 1306 1733 1326
rect 1682 1303 1701 1306
rect 1698 1216 1701 1303
rect 1722 1303 1733 1306
rect 1698 1213 1717 1216
rect 1642 1193 1645 1206
rect 1650 1166 1653 1206
rect 1642 1163 1653 1166
rect 1626 1133 1629 1156
rect 1610 1063 1621 1066
rect 1610 1013 1613 1056
rect 1570 1003 1581 1006
rect 1586 1003 1605 1006
rect 1610 983 1613 1006
rect 1514 973 1525 976
rect 1442 813 1445 846
rect 1450 826 1453 933
rect 1458 923 1469 926
rect 1474 853 1477 926
rect 1450 823 1461 826
rect 1474 813 1477 836
rect 1482 813 1485 926
rect 1490 913 1493 936
rect 1498 903 1501 926
rect 1506 813 1509 956
rect 1522 933 1525 973
rect 1618 963 1621 1063
rect 1626 953 1629 1126
rect 1634 1103 1637 1136
rect 1642 1113 1645 1163
rect 1698 1153 1701 1206
rect 1706 1183 1709 1206
rect 1714 1153 1717 1213
rect 1722 1183 1725 1303
rect 1762 1273 1765 1326
rect 1786 1236 1789 1326
rect 1794 1323 1797 1336
rect 1842 1333 1861 1336
rect 1818 1293 1821 1326
rect 1850 1313 1853 1333
rect 1858 1303 1861 1326
rect 1786 1233 1797 1236
rect 1746 1213 1749 1226
rect 1786 1213 1789 1226
rect 1730 1186 1733 1206
rect 1730 1183 1749 1186
rect 1730 1153 1733 1176
rect 1690 1133 1693 1146
rect 1674 1113 1677 1126
rect 1634 1013 1637 1026
rect 1682 1013 1685 1026
rect 1634 993 1637 1006
rect 1514 866 1517 926
rect 1522 913 1525 926
rect 1514 863 1525 866
rect 1530 853 1533 936
rect 1538 883 1541 926
rect 1546 916 1549 936
rect 1554 933 1557 946
rect 1554 923 1565 926
rect 1570 923 1573 936
rect 1546 913 1557 916
rect 1578 893 1581 926
rect 1586 883 1589 936
rect 1594 933 1597 946
rect 1650 933 1653 946
rect 1602 906 1605 926
rect 1626 923 1637 926
rect 1594 876 1597 906
rect 1602 903 1613 906
rect 1442 733 1445 786
rect 1474 763 1477 806
rect 1482 753 1485 806
rect 1490 763 1493 786
rect 1522 766 1525 786
rect 1506 763 1525 766
rect 1450 733 1453 746
rect 1442 663 1445 726
rect 1402 613 1405 656
rect 1426 613 1429 626
rect 1450 613 1453 726
rect 1474 673 1477 726
rect 1394 603 1405 606
rect 1394 596 1397 603
rect 1378 593 1397 596
rect 1402 583 1405 603
rect 1450 586 1453 606
rect 1426 583 1453 586
rect 1354 543 1373 546
rect 1354 533 1357 543
rect 1362 476 1365 536
rect 1370 533 1373 543
rect 1378 523 1381 546
rect 1426 533 1429 583
rect 1434 533 1437 566
rect 1458 553 1461 606
rect 1466 573 1469 626
rect 1474 603 1477 616
rect 1482 603 1485 636
rect 1498 613 1501 736
rect 1506 733 1509 763
rect 1514 733 1517 756
rect 1522 733 1525 746
rect 1530 733 1533 806
rect 1538 783 1541 876
rect 1586 873 1597 876
rect 1562 813 1565 856
rect 1570 813 1573 836
rect 1506 713 1509 726
rect 1514 676 1517 706
rect 1522 686 1525 726
rect 1530 713 1533 726
rect 1522 683 1533 686
rect 1514 673 1525 676
rect 1506 613 1509 626
rect 1514 606 1517 666
rect 1490 583 1493 606
rect 1498 603 1517 606
rect 1522 603 1525 673
rect 1530 613 1533 683
rect 1538 613 1541 756
rect 1554 733 1557 746
rect 1546 713 1549 726
rect 1562 713 1565 726
rect 1570 693 1573 786
rect 1578 703 1581 736
rect 1498 536 1501 596
rect 1394 513 1397 526
rect 1354 473 1365 476
rect 1346 423 1349 446
rect 1338 413 1349 416
rect 1354 413 1357 473
rect 1394 436 1397 506
rect 1386 433 1397 436
rect 1402 433 1405 526
rect 1370 413 1373 426
rect 1386 423 1389 433
rect 1194 333 1213 336
rect 1186 313 1189 326
rect 1202 276 1205 326
rect 1210 316 1213 333
rect 1218 323 1221 396
rect 1226 393 1237 396
rect 1226 333 1229 393
rect 1226 316 1229 326
rect 1210 313 1229 316
rect 1174 233 1181 236
rect 1178 216 1181 233
rect 1146 213 1157 216
rect 1162 183 1165 216
rect 1170 213 1181 216
rect 1186 213 1189 276
rect 1202 273 1213 276
rect 1170 156 1173 213
rect 1194 206 1197 256
rect 1178 176 1181 206
rect 1186 203 1197 206
rect 1202 206 1205 266
rect 1210 213 1213 273
rect 1218 216 1221 296
rect 1234 273 1237 336
rect 1242 266 1245 326
rect 1226 263 1245 266
rect 1226 223 1229 263
rect 1218 213 1229 216
rect 1234 213 1237 226
rect 1202 203 1213 206
rect 1186 186 1189 203
rect 1186 183 1197 186
rect 1178 173 1189 176
rect 1170 153 1181 156
rect 1178 133 1181 153
rect 1186 133 1189 173
rect 1146 53 1149 126
rect 1178 113 1181 126
rect 1186 103 1189 126
rect 1194 93 1197 183
rect 1202 143 1205 186
rect 1210 133 1213 203
rect 1218 133 1221 206
rect 1202 83 1205 126
rect 1210 93 1213 126
rect 1218 113 1221 126
rect 1226 106 1229 213
rect 1242 173 1245 236
rect 1250 223 1253 366
rect 1258 323 1261 346
rect 1258 203 1261 306
rect 1266 293 1269 376
rect 1274 263 1277 366
rect 1282 333 1285 396
rect 1322 356 1325 413
rect 1330 403 1341 406
rect 1322 353 1333 356
rect 1274 213 1277 226
rect 1266 173 1269 206
rect 1282 183 1285 276
rect 1242 156 1245 166
rect 1242 153 1277 156
rect 1274 133 1277 153
rect 1290 133 1293 216
rect 1298 213 1301 276
rect 1330 233 1333 353
rect 1338 313 1341 403
rect 1346 396 1349 413
rect 1346 393 1353 396
rect 1350 306 1353 393
rect 1402 363 1405 426
rect 1410 423 1413 446
rect 1418 433 1421 496
rect 1346 303 1353 306
rect 1362 303 1365 326
rect 1370 323 1373 336
rect 1378 333 1381 356
rect 1386 333 1397 336
rect 1386 316 1389 333
rect 1382 313 1389 316
rect 1346 253 1349 303
rect 1382 246 1385 313
rect 1394 303 1397 316
rect 1402 296 1405 346
rect 1410 333 1413 346
rect 1426 336 1429 516
rect 1434 493 1437 526
rect 1458 483 1461 526
rect 1466 473 1469 526
rect 1482 456 1485 536
rect 1490 533 1509 536
rect 1506 503 1509 526
rect 1514 523 1517 536
rect 1522 523 1525 596
rect 1538 583 1541 606
rect 1546 576 1549 636
rect 1554 613 1557 626
rect 1578 613 1581 636
rect 1586 613 1589 873
rect 1602 836 1605 896
rect 1594 833 1605 836
rect 1594 803 1597 833
rect 1610 816 1613 903
rect 1650 866 1653 926
rect 1658 903 1661 936
rect 1666 876 1669 926
rect 1674 903 1677 986
rect 1682 953 1685 1006
rect 1682 923 1685 946
rect 1690 933 1693 1126
rect 1698 1043 1701 1136
rect 1730 1046 1733 1126
rect 1746 1113 1749 1183
rect 1762 1133 1765 1146
rect 1730 1043 1741 1046
rect 1706 1013 1709 1026
rect 1738 993 1741 1043
rect 1754 1013 1757 1126
rect 1762 1013 1765 1126
rect 1770 1123 1773 1186
rect 1778 1103 1781 1206
rect 1794 1203 1797 1233
rect 1802 1183 1805 1196
rect 1810 1153 1813 1226
rect 1866 1213 1869 1416
rect 1906 1413 1909 1446
rect 1882 1333 1885 1346
rect 1882 1213 1885 1236
rect 1890 1213 1893 1336
rect 1914 1323 1917 1336
rect 1938 1333 1941 1406
rect 1922 1223 1925 1326
rect 1786 1113 1789 1126
rect 1658 873 1669 876
rect 1690 866 1693 926
rect 1714 903 1717 926
rect 1650 863 1669 866
rect 1610 813 1621 816
rect 1642 813 1645 826
rect 1650 813 1661 816
rect 1666 813 1669 863
rect 1674 863 1693 866
rect 1594 733 1597 796
rect 1642 773 1645 806
rect 1618 736 1621 746
rect 1618 733 1645 736
rect 1602 723 1613 726
rect 1618 716 1621 726
rect 1594 713 1621 716
rect 1626 713 1629 726
rect 1642 723 1645 733
rect 1642 673 1645 716
rect 1650 643 1653 806
rect 1658 793 1661 813
rect 1666 753 1669 806
rect 1674 763 1677 863
rect 1682 793 1685 806
rect 1690 756 1693 826
rect 1714 813 1717 866
rect 1722 813 1725 926
rect 1738 823 1741 936
rect 1746 866 1749 1006
rect 1754 953 1757 1006
rect 1770 993 1773 1036
rect 1778 1013 1781 1026
rect 1786 956 1789 1076
rect 1794 1063 1797 1136
rect 1842 1133 1845 1156
rect 1858 1146 1861 1206
rect 1866 1156 1869 1206
rect 1866 1153 1885 1156
rect 1858 1143 1869 1146
rect 1842 1113 1845 1126
rect 1850 1056 1853 1136
rect 1858 1106 1861 1136
rect 1866 1123 1869 1143
rect 1858 1103 1865 1106
rect 1842 1053 1853 1056
rect 1834 1003 1837 1016
rect 1842 1013 1845 1053
rect 1862 1036 1865 1103
rect 1874 1083 1877 1146
rect 1882 1113 1885 1153
rect 1890 1143 1893 1186
rect 1914 1163 1917 1206
rect 1922 1153 1925 1216
rect 1938 1213 1941 1316
rect 1946 1306 1949 1326
rect 1946 1303 1953 1306
rect 1950 1226 1953 1303
rect 1946 1223 1953 1226
rect 1946 1146 1949 1223
rect 1946 1143 1953 1146
rect 1858 1033 1865 1036
rect 1858 1013 1861 1033
rect 1890 1013 1893 1136
rect 1906 1113 1909 1126
rect 1842 956 1845 1006
rect 1890 983 1893 1006
rect 1786 953 1797 956
rect 1794 943 1797 953
rect 1802 936 1805 956
rect 1842 953 1853 956
rect 1794 933 1805 936
rect 1770 913 1773 926
rect 1754 873 1765 876
rect 1746 863 1757 866
rect 1690 753 1701 756
rect 1698 733 1701 753
rect 1706 733 1709 786
rect 1738 763 1741 816
rect 1746 813 1749 856
rect 1746 753 1749 806
rect 1754 803 1757 863
rect 1762 823 1765 873
rect 1762 796 1765 816
rect 1770 803 1773 876
rect 1778 813 1781 926
rect 1794 906 1797 926
rect 1786 903 1797 906
rect 1786 813 1789 903
rect 1802 866 1805 926
rect 1834 883 1837 926
rect 1802 863 1813 866
rect 1850 863 1853 953
rect 1778 796 1781 806
rect 1762 793 1781 796
rect 1762 783 1781 786
rect 1762 733 1765 783
rect 1794 763 1797 826
rect 1802 756 1805 836
rect 1810 803 1813 863
rect 1818 843 1837 846
rect 1818 823 1821 843
rect 1834 823 1837 843
rect 1850 833 1853 846
rect 1858 833 1861 976
rect 1818 796 1821 806
rect 1810 793 1821 796
rect 1826 793 1829 816
rect 1842 806 1845 826
rect 1866 823 1869 946
rect 1874 933 1877 956
rect 1882 933 1885 946
rect 1890 933 1893 966
rect 1898 953 1901 1096
rect 1906 973 1909 1056
rect 1914 1013 1917 1026
rect 1922 1003 1925 1106
rect 1938 1096 1941 1136
rect 1930 1093 1941 1096
rect 1930 1053 1933 1093
rect 1930 993 1933 1016
rect 1914 953 1917 986
rect 1938 943 1941 1086
rect 1950 1046 1953 1143
rect 1946 1043 1953 1046
rect 1946 1023 1949 1043
rect 1946 986 1949 1006
rect 1946 983 1953 986
rect 1874 843 1877 926
rect 1834 803 1845 806
rect 1794 753 1805 756
rect 1810 733 1813 756
rect 1818 733 1821 793
rect 1602 603 1605 626
rect 1538 573 1549 576
rect 1610 573 1613 606
rect 1658 603 1661 706
rect 1674 696 1677 726
rect 1666 693 1677 696
rect 1666 613 1677 616
rect 1682 613 1685 726
rect 1666 596 1669 606
rect 1658 593 1669 596
rect 1474 453 1485 456
rect 1434 393 1437 426
rect 1442 413 1461 416
rect 1418 333 1429 336
rect 1434 333 1437 366
rect 1442 353 1445 413
rect 1450 403 1461 406
rect 1450 376 1453 403
rect 1450 373 1461 376
rect 1466 373 1469 436
rect 1442 333 1445 346
rect 1418 303 1421 333
rect 1394 293 1405 296
rect 1382 243 1389 246
rect 1306 213 1317 216
rect 1298 163 1301 206
rect 1306 203 1317 206
rect 1218 103 1229 106
rect 1250 103 1253 126
rect 1282 113 1285 126
rect 1298 123 1301 136
rect 1306 133 1309 203
rect 1322 193 1325 206
rect 1314 133 1317 176
rect 1330 173 1333 216
rect 1338 213 1341 226
rect 1362 213 1365 226
rect 1386 213 1389 243
rect 1338 193 1341 206
rect 1186 0 1189 46
rect 1202 0 1205 26
rect 1218 0 1221 103
rect 1250 0 1253 66
rect 1266 0 1269 96
rect 1314 93 1317 126
rect 1322 103 1325 126
rect 1346 113 1349 126
rect 1378 123 1381 176
rect 1386 103 1389 126
rect 1282 0 1285 56
rect 1362 0 1365 16
rect 1394 13 1397 293
rect 1418 213 1421 226
rect 1426 213 1429 326
rect 1434 256 1437 326
rect 1434 253 1445 256
rect 1442 213 1445 253
rect 1450 233 1453 336
rect 1458 243 1461 373
rect 1466 333 1469 356
rect 1474 333 1477 453
rect 1482 393 1485 416
rect 1490 403 1493 496
rect 1498 363 1501 416
rect 1506 353 1509 426
rect 1514 413 1517 496
rect 1522 413 1525 476
rect 1530 433 1533 536
rect 1538 503 1541 573
rect 1546 456 1549 526
rect 1570 516 1573 526
rect 1562 513 1573 516
rect 1562 483 1565 513
rect 1546 453 1557 456
rect 1554 413 1557 453
rect 1570 413 1573 506
rect 1578 493 1581 526
rect 1594 513 1597 536
rect 1602 533 1605 546
rect 1650 533 1653 566
rect 1658 526 1661 593
rect 1674 586 1677 613
rect 1690 603 1693 676
rect 1698 613 1701 726
rect 1706 693 1709 726
rect 1730 703 1733 726
rect 1738 713 1741 726
rect 1730 613 1733 666
rect 1754 613 1757 726
rect 1786 713 1789 726
rect 1514 403 1525 406
rect 1522 333 1525 403
rect 1530 333 1533 376
rect 1474 313 1477 326
rect 1498 313 1501 326
rect 1554 323 1565 326
rect 1450 216 1453 226
rect 1450 213 1461 216
rect 1450 193 1453 206
rect 1402 113 1405 126
rect 1410 113 1413 126
rect 1402 103 1413 106
rect 1418 103 1421 126
rect 1426 123 1429 166
rect 1434 113 1437 176
rect 1458 173 1461 213
rect 1466 153 1469 216
rect 1474 173 1477 206
rect 1482 203 1485 236
rect 1530 213 1533 316
rect 1578 286 1581 416
rect 1602 413 1605 526
rect 1650 523 1661 526
rect 1650 413 1653 523
rect 1666 506 1669 586
rect 1674 583 1685 586
rect 1682 533 1685 583
rect 1662 503 1669 506
rect 1662 436 1665 503
rect 1662 433 1669 436
rect 1674 433 1677 526
rect 1690 483 1693 596
rect 1698 533 1701 606
rect 1706 553 1709 606
rect 1754 586 1757 606
rect 1762 603 1765 646
rect 1778 643 1781 706
rect 1794 673 1797 726
rect 1810 653 1813 726
rect 1826 723 1829 766
rect 1834 726 1837 803
rect 1842 733 1845 786
rect 1850 773 1853 816
rect 1858 793 1861 816
rect 1834 723 1845 726
rect 1818 613 1821 626
rect 1746 583 1757 586
rect 1722 483 1725 526
rect 1666 413 1669 433
rect 1586 403 1597 406
rect 1586 333 1589 396
rect 1634 333 1637 376
rect 1642 343 1645 356
rect 1650 343 1653 406
rect 1658 373 1661 406
rect 1666 393 1669 406
rect 1578 283 1589 286
rect 1538 206 1541 216
rect 1554 213 1557 226
rect 1586 213 1589 283
rect 1610 223 1613 326
rect 1618 213 1621 276
rect 1642 213 1645 336
rect 1650 333 1661 336
rect 1666 323 1669 356
rect 1674 346 1677 416
rect 1682 403 1685 476
rect 1690 413 1693 426
rect 1698 353 1701 436
rect 1674 343 1685 346
rect 1674 313 1677 336
rect 1674 226 1677 246
rect 1650 223 1677 226
rect 1658 213 1669 216
rect 1674 213 1677 223
rect 1682 206 1685 343
rect 1690 333 1693 346
rect 1698 213 1701 326
rect 1706 233 1709 446
rect 1746 433 1749 583
rect 1762 543 1765 596
rect 1754 533 1765 536
rect 1770 533 1773 586
rect 1810 556 1813 606
rect 1818 573 1821 606
rect 1826 566 1829 716
rect 1842 713 1845 723
rect 1834 593 1837 696
rect 1842 583 1845 656
rect 1850 613 1853 736
rect 1858 733 1861 746
rect 1866 726 1869 776
rect 1874 763 1877 816
rect 1882 756 1885 806
rect 1890 773 1893 926
rect 1914 913 1917 926
rect 1906 823 1909 906
rect 1922 813 1925 926
rect 1938 816 1941 936
rect 1950 826 1953 983
rect 1950 823 1957 826
rect 1938 813 1949 816
rect 1858 723 1869 726
rect 1874 753 1885 756
rect 1874 723 1877 753
rect 1882 733 1885 746
rect 1890 733 1893 756
rect 1898 733 1901 746
rect 1858 713 1861 723
rect 1858 603 1861 616
rect 1866 613 1869 626
rect 1778 553 1813 556
rect 1818 563 1829 566
rect 1834 563 1861 566
rect 1874 563 1877 716
rect 1906 706 1909 776
rect 1930 746 1933 786
rect 1938 773 1941 806
rect 1898 703 1909 706
rect 1898 646 1901 703
rect 1898 643 1909 646
rect 1882 573 1885 626
rect 1906 613 1909 643
rect 1914 623 1917 736
rect 1922 723 1925 746
rect 1930 743 1941 746
rect 1930 713 1933 736
rect 1938 686 1941 743
rect 1946 723 1949 813
rect 1954 706 1957 823
rect 1946 703 1957 706
rect 1946 693 1949 703
rect 1930 683 1941 686
rect 1930 663 1933 683
rect 1930 613 1933 646
rect 1930 573 1933 596
rect 1754 493 1757 533
rect 1730 413 1741 416
rect 1754 413 1757 486
rect 1762 443 1765 526
rect 1770 473 1773 526
rect 1762 413 1765 436
rect 1778 423 1781 553
rect 1786 513 1789 526
rect 1794 506 1797 536
rect 1802 533 1813 536
rect 1818 533 1821 563
rect 1834 556 1837 563
rect 1826 553 1837 556
rect 1858 556 1861 563
rect 1858 553 1877 556
rect 1826 533 1829 553
rect 1874 533 1877 553
rect 1802 523 1813 526
rect 1786 503 1797 506
rect 1786 433 1789 503
rect 1794 413 1797 496
rect 1714 206 1717 386
rect 1722 316 1725 366
rect 1722 313 1729 316
rect 1738 313 1741 326
rect 1726 246 1729 313
rect 1746 263 1749 356
rect 1754 333 1757 406
rect 1762 386 1765 406
rect 1810 403 1813 516
rect 1818 503 1821 526
rect 1826 513 1829 526
rect 1818 396 1821 406
rect 1826 403 1829 476
rect 1882 466 1885 536
rect 1882 463 1893 466
rect 1834 403 1837 416
rect 1882 413 1885 456
rect 1890 413 1893 463
rect 1898 436 1901 526
rect 1914 443 1917 516
rect 1898 433 1909 436
rect 1762 383 1773 386
rect 1762 293 1765 376
rect 1770 306 1773 383
rect 1778 333 1781 386
rect 1810 353 1813 396
rect 1818 393 1829 396
rect 1842 393 1845 406
rect 1826 333 1829 393
rect 1850 383 1853 406
rect 1858 356 1861 406
rect 1858 353 1885 356
rect 1834 333 1837 346
rect 1810 306 1813 326
rect 1834 313 1837 326
rect 1770 303 1789 306
rect 1810 303 1821 306
rect 1858 303 1861 326
rect 1882 316 1885 353
rect 1890 323 1893 386
rect 1906 353 1909 433
rect 1930 413 1933 526
rect 1914 393 1917 406
rect 1882 313 1893 316
rect 1722 243 1729 246
rect 1722 223 1725 243
rect 1730 216 1733 226
rect 1530 203 1541 206
rect 1594 193 1597 206
rect 1442 113 1445 136
rect 1458 113 1461 126
rect 1514 123 1517 156
rect 1522 136 1525 176
rect 1522 133 1533 136
rect 1498 103 1501 116
rect 1522 83 1525 133
rect 1530 103 1533 126
rect 1546 113 1549 156
rect 1602 133 1605 166
rect 1650 163 1653 206
rect 1674 196 1677 206
rect 1682 203 1701 206
rect 1706 203 1717 206
rect 1722 213 1733 216
rect 1738 213 1741 236
rect 1754 213 1765 216
rect 1786 213 1789 303
rect 1794 213 1797 226
rect 1818 213 1821 303
rect 1674 193 1685 196
rect 1554 113 1557 126
rect 1570 123 1581 126
rect 1610 103 1613 126
rect 1634 93 1637 126
rect 1642 113 1645 126
rect 1658 123 1661 136
rect 1666 113 1669 186
rect 1682 106 1685 193
rect 1706 173 1709 203
rect 1722 196 1725 213
rect 1714 193 1725 196
rect 1730 193 1733 206
rect 1690 113 1693 136
rect 1706 123 1709 166
rect 1714 116 1717 193
rect 1730 133 1733 176
rect 1746 153 1749 186
rect 1778 133 1781 146
rect 1722 123 1733 126
rect 1714 113 1725 116
rect 1682 103 1693 106
rect 1786 73 1789 206
rect 1794 163 1797 206
rect 1794 133 1797 146
rect 1810 133 1813 186
rect 1842 183 1845 296
rect 1858 213 1861 266
rect 1882 236 1885 306
rect 1866 233 1885 236
rect 1866 223 1869 233
rect 1850 203 1869 206
rect 1818 126 1821 176
rect 1850 173 1853 203
rect 1802 123 1821 126
rect 1826 123 1829 166
rect 1834 123 1837 156
rect 1850 113 1853 166
rect 1858 143 1861 196
rect 1874 163 1877 226
rect 1882 153 1885 233
rect 1890 206 1893 313
rect 1898 213 1901 226
rect 1890 203 1901 206
rect 1906 196 1909 326
rect 1938 283 1941 676
rect 1946 603 1949 616
rect 1946 556 1949 576
rect 1946 553 1953 556
rect 1950 386 1953 553
rect 1946 383 1953 386
rect 1946 363 1949 383
rect 1914 233 1917 256
rect 1914 213 1917 226
rect 1906 193 1917 196
rect 1914 133 1917 193
rect 1890 113 1893 126
rect 1906 123 1917 126
rect 1922 123 1925 236
rect 1930 213 1933 226
rect 1930 123 1941 126
rect 1960 37 1980 1903
rect 1984 13 2004 1927
rect 2010 946 2013 966
rect 2010 943 2017 946
rect 2014 756 2017 943
rect 2010 753 2017 756
rect 2010 733 2013 753
rect 2010 706 2013 726
rect 2010 703 2017 706
rect 2014 566 2017 703
rect 2010 563 2017 566
rect 2010 543 2013 563
rect 2010 493 2013 536
<< metal3 >>
rect 1297 1922 1326 1927
rect 1329 1912 1398 1917
rect 969 1902 1070 1907
rect 1393 1902 1526 1907
rect 953 1892 1054 1897
rect 937 1882 1086 1887
rect 761 1872 846 1877
rect 905 1872 1022 1877
rect 1441 1872 1574 1877
rect 825 1862 902 1867
rect 921 1862 1046 1867
rect 1273 1862 1398 1867
rect 1273 1857 1278 1862
rect 769 1852 870 1857
rect 889 1852 1038 1857
rect 1249 1852 1278 1857
rect 1393 1857 1398 1862
rect 1441 1857 1446 1872
rect 1393 1852 1446 1857
rect 1569 1857 1574 1872
rect 1569 1852 1822 1857
rect 729 1842 974 1847
rect 1201 1842 1342 1847
rect 1425 1842 1558 1847
rect 1201 1837 1206 1842
rect 177 1832 214 1837
rect 657 1832 694 1837
rect 737 1832 790 1837
rect 833 1832 894 1837
rect 953 1832 1206 1837
rect 1217 1832 1278 1837
rect 1369 1832 1510 1837
rect 289 1822 342 1827
rect 609 1822 678 1827
rect 801 1822 862 1827
rect 873 1822 966 1827
rect 977 1822 1030 1827
rect 1177 1822 1230 1827
rect 1385 1822 1430 1827
rect 1441 1822 1486 1827
rect 1577 1822 1646 1827
rect 1689 1822 1742 1827
rect 1833 1822 1942 1827
rect 0 1812 174 1817
rect 577 1812 774 1817
rect 257 1802 310 1807
rect 385 1802 486 1807
rect 505 1802 534 1807
rect 545 1802 582 1807
rect 601 1802 718 1807
rect 801 1802 806 1822
rect 1577 1817 1582 1822
rect 913 1812 1006 1817
rect 1297 1812 1350 1817
rect 1401 1812 1582 1817
rect 1641 1817 1646 1822
rect 1641 1812 1806 1817
rect 977 1802 1070 1807
rect 1249 1802 1366 1807
rect 1481 1802 1534 1807
rect 1593 1802 1646 1807
rect 1697 1802 1750 1807
rect 385 1797 390 1802
rect 129 1792 214 1797
rect 361 1792 390 1797
rect 481 1797 486 1802
rect 1249 1797 1254 1802
rect 1361 1797 1366 1802
rect 481 1792 558 1797
rect 585 1792 614 1797
rect 641 1792 758 1797
rect 849 1792 942 1797
rect 1113 1792 1254 1797
rect 1273 1792 1350 1797
rect 1361 1792 1462 1797
rect 1553 1792 1582 1797
rect 1577 1787 1582 1792
rect 1753 1792 1862 1797
rect 1753 1787 1758 1792
rect 281 1782 406 1787
rect 681 1782 742 1787
rect 753 1782 990 1787
rect 1265 1782 1398 1787
rect 1577 1782 1758 1787
rect 321 1772 478 1777
rect 561 1772 590 1777
rect 793 1772 870 1777
rect 1777 1772 1870 1777
rect 609 1767 702 1772
rect 889 1767 1014 1772
rect 305 1762 334 1767
rect 385 1762 446 1767
rect 473 1762 614 1767
rect 697 1762 894 1767
rect 1009 1762 1038 1767
rect 1273 1762 1326 1767
rect 1521 1762 1734 1767
rect 1521 1757 1526 1762
rect 233 1752 302 1757
rect 401 1752 614 1757
rect 641 1752 686 1757
rect 761 1752 798 1757
rect 809 1752 838 1757
rect 857 1752 1134 1757
rect 1353 1752 1526 1757
rect 1729 1757 1734 1762
rect 1729 1752 1758 1757
rect 129 1742 190 1747
rect 249 1742 430 1747
rect 481 1742 558 1747
rect 577 1742 622 1747
rect 665 1742 726 1747
rect 785 1742 838 1747
rect 969 1742 1006 1747
rect 1089 1742 1390 1747
rect 1585 1742 1654 1747
rect 1585 1737 1590 1742
rect 0 1732 182 1737
rect 417 1732 494 1737
rect 625 1732 662 1737
rect 673 1732 726 1737
rect 881 1732 918 1737
rect 1033 1732 1078 1737
rect 1537 1732 1590 1737
rect 1649 1737 1654 1742
rect 1649 1732 1718 1737
rect 265 1722 302 1727
rect 505 1722 534 1727
rect 857 1722 878 1727
rect 1065 1722 1118 1727
rect 1601 1722 1638 1727
rect 321 1712 406 1717
rect 513 1712 582 1717
rect 681 1712 766 1717
rect 857 1712 886 1717
rect 1017 1712 1078 1717
rect 1193 1712 1246 1717
rect 1369 1712 1438 1717
rect 1457 1712 1502 1717
rect 1785 1712 1870 1717
rect 1369 1707 1374 1712
rect 185 1702 238 1707
rect 353 1702 486 1707
rect 521 1702 574 1707
rect 641 1702 742 1707
rect 1137 1702 1262 1707
rect 1345 1702 1374 1707
rect 1433 1707 1438 1712
rect 1433 1702 1494 1707
rect 225 1692 294 1697
rect 417 1692 534 1697
rect 609 1692 662 1697
rect 721 1692 966 1697
rect 1345 1692 1454 1697
rect 561 1682 590 1687
rect 1257 1682 1414 1687
rect 1409 1677 1414 1682
rect 1505 1682 1902 1687
rect 1505 1677 1510 1682
rect 1409 1672 1510 1677
rect 1745 1672 1774 1677
rect 1769 1667 1774 1672
rect 1865 1672 1894 1677
rect 1865 1667 1870 1672
rect 753 1662 1014 1667
rect 1769 1662 1870 1667
rect 249 1652 286 1657
rect 449 1652 710 1657
rect 449 1637 454 1652
rect 265 1632 358 1637
rect 425 1632 454 1637
rect 705 1637 710 1652
rect 753 1647 758 1662
rect 729 1642 758 1647
rect 1009 1647 1014 1662
rect 1177 1652 1390 1657
rect 1009 1642 1070 1647
rect 705 1632 742 1637
rect 801 1632 854 1637
rect 897 1632 1030 1637
rect 1281 1632 1318 1637
rect 353 1627 358 1632
rect 129 1622 174 1627
rect 353 1622 422 1627
rect 465 1622 510 1627
rect 625 1622 678 1627
rect 697 1622 806 1627
rect 833 1622 870 1627
rect 1017 1622 1054 1627
rect 1105 1622 1158 1627
rect 417 1617 422 1622
rect 177 1612 230 1617
rect 249 1612 310 1617
rect 345 1612 406 1617
rect 417 1612 486 1617
rect 713 1612 742 1617
rect 225 1607 230 1612
rect 225 1602 326 1607
rect 505 1602 694 1607
rect 737 1602 742 1612
rect 945 1607 950 1617
rect 985 1612 1046 1617
rect 1249 1612 1294 1617
rect 785 1602 878 1607
rect 897 1602 950 1607
rect 1001 1602 1094 1607
rect 1161 1602 1278 1607
rect 505 1597 510 1602
rect 153 1592 270 1597
rect 441 1592 510 1597
rect 689 1597 694 1602
rect 785 1597 790 1602
rect 689 1592 790 1597
rect 873 1597 878 1602
rect 1313 1597 1318 1627
rect 1337 1622 1422 1627
rect 1561 1622 1614 1627
rect 1705 1622 1758 1627
rect 1393 1602 1470 1607
rect 1761 1602 1854 1607
rect 1969 1602 2020 1607
rect 1761 1597 1766 1602
rect 1969 1597 1974 1602
rect 873 1592 1102 1597
rect 1313 1592 1342 1597
rect 1497 1592 1566 1597
rect 1617 1592 1766 1597
rect 1777 1592 1974 1597
rect 529 1587 670 1592
rect 481 1582 534 1587
rect 665 1582 734 1587
rect 801 1582 902 1587
rect 929 1582 966 1587
rect 1009 1582 1038 1587
rect 1409 1582 1462 1587
rect 1521 1582 1670 1587
rect 457 1572 934 1577
rect 1049 1572 1430 1577
rect 929 1567 1054 1572
rect 1425 1567 1430 1572
rect 1537 1572 1798 1577
rect 1537 1567 1542 1572
rect 657 1562 910 1567
rect 1425 1562 1542 1567
rect 1561 1562 1670 1567
rect 561 1557 638 1562
rect 1201 1557 1270 1562
rect 1665 1557 1670 1562
rect 1753 1562 1862 1567
rect 1753 1557 1758 1562
rect 89 1552 238 1557
rect 385 1552 446 1557
rect 481 1552 566 1557
rect 633 1552 822 1557
rect 953 1552 1206 1557
rect 1265 1552 1382 1557
rect 1601 1552 1630 1557
rect 1665 1552 1758 1557
rect 89 1537 94 1552
rect 65 1532 94 1537
rect 233 1537 238 1552
rect 257 1542 286 1547
rect 305 1542 342 1547
rect 425 1542 470 1547
rect 577 1542 686 1547
rect 745 1542 838 1547
rect 1217 1542 1334 1547
rect 1377 1542 1646 1547
rect 233 1532 382 1537
rect 713 1532 742 1537
rect 993 1532 1054 1537
rect 1097 1532 1206 1537
rect 1745 1532 1790 1537
rect 65 1527 70 1532
rect 0 1522 70 1527
rect 81 1522 158 1527
rect 281 1522 334 1527
rect 345 1522 390 1527
rect 1017 1522 1046 1527
rect 1601 1522 1758 1527
rect 217 1512 294 1517
rect 353 1512 478 1517
rect 553 1512 622 1517
rect 729 1512 782 1517
rect 929 1512 958 1517
rect 1105 1512 1150 1517
rect 1265 1512 1310 1517
rect 1361 1512 1406 1517
rect 1537 1512 1582 1517
rect 1753 1512 1814 1517
rect 1841 1512 1886 1517
rect 1905 1512 2020 1517
rect 1905 1507 1910 1512
rect 313 1502 374 1507
rect 393 1502 422 1507
rect 417 1497 422 1502
rect 489 1502 534 1507
rect 561 1502 686 1507
rect 825 1502 982 1507
rect 1025 1502 1126 1507
rect 1481 1502 1590 1507
rect 1849 1502 1910 1507
rect 489 1497 494 1502
rect 337 1492 358 1497
rect 417 1492 494 1497
rect 521 1492 550 1497
rect 545 1487 550 1492
rect 617 1492 726 1497
rect 617 1487 622 1492
rect 201 1482 286 1487
rect 545 1482 622 1487
rect 0 1472 318 1477
rect 1009 1472 1086 1477
rect 481 1462 678 1467
rect 217 1452 278 1457
rect 481 1447 486 1462
rect 337 1442 446 1447
rect 457 1442 486 1447
rect 673 1447 678 1462
rect 841 1462 950 1467
rect 841 1457 846 1462
rect 817 1452 846 1457
rect 945 1457 950 1462
rect 945 1452 1038 1457
rect 1585 1452 1870 1457
rect 1585 1447 1590 1452
rect 673 1442 702 1447
rect 1257 1442 1326 1447
rect 1561 1442 1590 1447
rect 1865 1447 1870 1452
rect 1865 1442 1910 1447
rect 1257 1437 1262 1442
rect 305 1432 382 1437
rect 473 1432 526 1437
rect 537 1432 574 1437
rect 657 1432 934 1437
rect 1193 1432 1262 1437
rect 1321 1437 1326 1442
rect 1321 1432 1350 1437
rect 1377 1432 1470 1437
rect 1761 1432 1854 1437
rect 369 1422 390 1427
rect 977 1422 1062 1427
rect 1273 1422 1302 1427
rect 1361 1422 1406 1427
rect 1505 1422 1534 1427
rect 1601 1422 1638 1427
rect 1649 1422 1718 1427
rect 1753 1422 1798 1427
rect 129 1412 222 1417
rect 321 1412 366 1417
rect 449 1412 550 1417
rect 1001 1412 1102 1417
rect 1505 1407 1510 1422
rect 1649 1417 1654 1422
rect 1585 1412 1654 1417
rect 385 1402 446 1407
rect 457 1402 486 1407
rect 569 1402 766 1407
rect 793 1402 846 1407
rect 913 1402 1054 1407
rect 1385 1402 1510 1407
rect 569 1397 574 1402
rect 425 1392 502 1397
rect 545 1392 574 1397
rect 761 1397 766 1402
rect 761 1392 838 1397
rect 849 1392 894 1397
rect 945 1392 990 1397
rect 1241 1392 1302 1397
rect 1329 1392 1374 1397
rect 1409 1392 1438 1397
rect 833 1387 838 1392
rect 1433 1387 1438 1392
rect 1521 1392 1582 1397
rect 1689 1392 1742 1397
rect 1521 1387 1526 1392
rect 337 1382 430 1387
rect 449 1382 622 1387
rect 641 1382 774 1387
rect 833 1382 998 1387
rect 449 1377 454 1382
rect 993 1377 998 1382
rect 1073 1382 1222 1387
rect 1377 1382 1398 1387
rect 1433 1382 1526 1387
rect 1601 1382 1646 1387
rect 1073 1377 1078 1382
rect 361 1372 454 1377
rect 545 1372 662 1377
rect 737 1372 942 1377
rect 993 1372 1078 1377
rect 1217 1377 1222 1382
rect 1217 1372 1358 1377
rect 113 1362 206 1367
rect 569 1362 830 1367
rect 1081 1362 1118 1367
rect 1129 1362 1150 1367
rect 1185 1362 1254 1367
rect 121 1352 230 1357
rect 473 1352 558 1357
rect 593 1352 750 1357
rect 809 1352 950 1357
rect 961 1352 1070 1357
rect 1201 1352 1246 1357
rect 25 1342 94 1347
rect 169 1342 302 1347
rect 25 1337 30 1342
rect 0 1332 30 1337
rect 89 1337 94 1342
rect 89 1332 294 1337
rect 561 1327 566 1347
rect 601 1342 654 1347
rect 681 1342 726 1347
rect 833 1342 870 1347
rect 937 1342 1022 1347
rect 657 1332 678 1337
rect 745 1332 806 1337
rect 89 1322 110 1327
rect 177 1322 254 1327
rect 273 1322 294 1327
rect 329 1322 358 1327
rect 545 1322 566 1327
rect 577 1322 638 1327
rect 673 1322 678 1332
rect 705 1322 766 1327
rect 817 1322 854 1327
rect 865 1317 870 1342
rect 1153 1337 1158 1347
rect 1169 1342 1270 1347
rect 1329 1337 1334 1372
rect 1417 1362 1550 1367
rect 1577 1362 1598 1367
rect 1417 1357 1422 1362
rect 1353 1352 1422 1357
rect 1545 1357 1550 1362
rect 1545 1352 1574 1357
rect 1777 1352 1862 1357
rect 1777 1347 1782 1352
rect 1345 1342 1414 1347
rect 1449 1342 1486 1347
rect 1513 1342 1550 1347
rect 1129 1332 1198 1337
rect 1329 1332 1350 1337
rect 1369 1332 1390 1337
rect 977 1322 1094 1327
rect 1137 1322 1238 1327
rect 0 1312 78 1317
rect 137 1312 166 1317
rect 185 1312 334 1317
rect 409 1312 430 1317
rect 561 1312 614 1317
rect 625 1312 662 1317
rect 681 1312 734 1317
rect 825 1312 870 1317
rect 1001 1312 1046 1317
rect 1385 1312 1390 1332
rect 1409 1312 1414 1342
rect 1665 1337 1670 1347
rect 1737 1342 1782 1347
rect 1857 1347 1862 1352
rect 1857 1342 1886 1347
rect 1473 1332 1534 1337
rect 73 1307 142 1312
rect 625 1307 630 1312
rect 1473 1307 1478 1332
rect 1553 1312 1558 1337
rect 1633 1332 1670 1337
rect 1857 1332 1894 1337
rect 1609 1322 1710 1327
rect 1793 1322 1870 1327
rect 1913 1322 1950 1327
rect 1593 1312 1630 1317
rect 169 1302 230 1307
rect 305 1302 462 1307
rect 569 1302 630 1307
rect 785 1302 854 1307
rect 1313 1302 1366 1307
rect 1473 1302 1590 1307
rect 1857 1302 1942 1307
rect 0 1292 182 1297
rect 249 1292 270 1297
rect 321 1292 366 1297
rect 385 1292 582 1297
rect 617 1292 718 1297
rect 729 1292 1390 1297
rect 1561 1292 1822 1297
rect 209 1282 430 1287
rect 537 1282 670 1287
rect 713 1282 830 1287
rect 1289 1282 1326 1287
rect 1537 1282 1582 1287
rect 0 1272 366 1277
rect 377 1272 598 1277
rect 761 1272 902 1277
rect 921 1272 1006 1277
rect 1105 1272 1134 1277
rect 1201 1272 1350 1277
rect 1409 1272 1494 1277
rect 1521 1272 1566 1277
rect 0 1252 5 1272
rect 921 1267 926 1272
rect 161 1262 390 1267
rect 417 1262 470 1267
rect 497 1262 646 1267
rect 657 1262 750 1267
rect 849 1262 926 1267
rect 1001 1267 1006 1272
rect 1409 1267 1414 1272
rect 1001 1262 1414 1267
rect 1489 1267 1494 1272
rect 1561 1267 1566 1272
rect 1737 1272 1766 1277
rect 1737 1267 1742 1272
rect 1489 1262 1518 1267
rect 1561 1262 1742 1267
rect 745 1257 854 1262
rect 337 1252 382 1257
rect 401 1252 558 1257
rect 657 1252 726 1257
rect 873 1252 990 1257
rect 1121 1252 1150 1257
rect 1257 1252 1326 1257
rect 1369 1252 1406 1257
rect 201 1247 318 1252
rect 1441 1247 1518 1252
rect 121 1242 206 1247
rect 313 1242 406 1247
rect 481 1242 878 1247
rect 1001 1242 1334 1247
rect 1417 1242 1446 1247
rect 1513 1242 1542 1247
rect 873 1237 1006 1242
rect 1329 1237 1422 1242
rect 217 1232 294 1237
rect 305 1232 550 1237
rect 601 1232 654 1237
rect 1097 1232 1126 1237
rect 1137 1232 1166 1237
rect 1457 1232 1510 1237
rect 1601 1232 1622 1237
rect 1881 1232 1926 1237
rect 729 1227 854 1232
rect 1201 1227 1310 1232
rect 0 1222 254 1227
rect 265 1222 302 1227
rect 329 1222 358 1227
rect 449 1222 502 1227
rect 529 1222 566 1227
rect 633 1222 694 1227
rect 705 1222 734 1227
rect 849 1222 878 1227
rect 905 1222 958 1227
rect 1001 1222 1046 1227
rect 1177 1222 1206 1227
rect 1305 1222 1334 1227
rect 1425 1222 1534 1227
rect 1673 1222 1750 1227
rect 1785 1222 1814 1227
rect 241 1212 318 1217
rect 345 1212 518 1217
rect 561 1212 806 1217
rect 825 1212 886 1217
rect 945 1212 966 1217
rect 977 1212 1094 1217
rect 1185 1212 1238 1217
rect 1281 1212 1382 1217
rect 1537 1212 1670 1217
rect 1865 1212 1926 1217
rect 1665 1207 1670 1212
rect 193 1202 230 1207
rect 377 1202 446 1207
rect 489 1202 550 1207
rect 817 1202 918 1207
rect 929 1202 1150 1207
rect 1201 1202 1310 1207
rect 1529 1202 1558 1207
rect 1665 1202 1830 1207
rect 1825 1197 1830 1202
rect 377 1192 462 1197
rect 617 1192 710 1197
rect 753 1192 1038 1197
rect 1169 1192 1246 1197
rect 1329 1192 1446 1197
rect 1513 1192 1550 1197
rect 1561 1192 1646 1197
rect 1825 1192 1878 1197
rect 1873 1187 1878 1192
rect 81 1182 158 1187
rect 225 1182 278 1187
rect 337 1182 374 1187
rect 433 1182 534 1187
rect 545 1182 630 1187
rect 745 1182 782 1187
rect 801 1182 998 1187
rect 1297 1182 1510 1187
rect 1609 1182 1710 1187
rect 1721 1182 1774 1187
rect 1801 1182 1862 1187
rect 1873 1182 1894 1187
rect 625 1177 726 1182
rect 0 1172 222 1177
rect 281 1172 422 1177
rect 457 1172 486 1177
rect 721 1172 942 1177
rect 993 1167 998 1182
rect 1009 1172 1054 1177
rect 1113 1172 1182 1177
rect 1201 1172 1390 1177
rect 1481 1172 1606 1177
rect 1697 1172 1734 1177
rect 1385 1167 1486 1172
rect 241 1162 502 1167
rect 553 1162 974 1167
rect 993 1162 1366 1167
rect 1505 1162 1782 1167
rect 1873 1162 1918 1167
rect 89 1157 182 1162
rect 0 1152 94 1157
rect 177 1152 230 1157
rect 249 1152 510 1157
rect 609 1152 1166 1157
rect 1193 1152 1270 1157
rect 1289 1152 1326 1157
rect 1465 1152 1502 1157
rect 1553 1152 1598 1157
rect 1625 1152 1702 1157
rect 129 1142 174 1147
rect 321 1142 342 1147
rect 409 1142 526 1147
rect 601 1142 686 1147
rect 697 1142 742 1147
rect 769 1142 814 1147
rect 865 1142 910 1147
rect 1129 1142 1214 1147
rect 1313 1142 1334 1147
rect 1345 1142 1382 1147
rect 1449 1142 1542 1147
rect 1601 1142 1694 1147
rect 929 1137 998 1142
rect 1041 1137 1110 1142
rect 1329 1137 1334 1142
rect 209 1132 390 1137
rect 425 1132 470 1137
rect 785 1132 806 1137
rect 849 1132 934 1137
rect 993 1132 1046 1137
rect 1105 1132 1142 1137
rect 1161 1132 1286 1137
rect 1329 1132 1518 1137
rect 1137 1127 1142 1132
rect 1281 1127 1286 1132
rect 1649 1127 1654 1142
rect 1713 1127 1718 1157
rect 121 1122 190 1127
rect 321 1122 358 1127
rect 505 1122 534 1127
rect 649 1122 822 1127
rect 833 1122 870 1127
rect 881 1122 982 1127
rect 1057 1122 1118 1127
rect 1137 1122 1190 1127
rect 1281 1122 1382 1127
rect 1625 1122 1654 1127
rect 1689 1122 1718 1127
rect 1729 1122 1734 1157
rect 1809 1152 1846 1157
rect 1873 1147 1878 1162
rect 1905 1152 1926 1157
rect 1761 1142 1878 1147
rect 1761 1132 1846 1137
rect 1761 1122 1766 1132
rect 1889 1127 1894 1147
rect 1857 1122 1894 1127
rect 817 1117 822 1122
rect 1401 1117 1510 1122
rect 273 1112 318 1117
rect 345 1112 414 1117
rect 481 1112 710 1117
rect 737 1112 806 1117
rect 817 1112 926 1117
rect 993 1112 1134 1117
rect 1145 1112 1182 1117
rect 1193 1112 1254 1117
rect 1305 1112 1406 1117
rect 1505 1112 1614 1117
rect 1641 1112 1678 1117
rect 1745 1112 1790 1117
rect 1841 1112 1886 1117
rect 1905 1112 1910 1152
rect 921 1107 998 1112
rect 217 1102 358 1107
rect 425 1102 462 1107
rect 521 1102 846 1107
rect 865 1102 902 1107
rect 1105 1102 1182 1107
rect 1193 1102 1246 1107
rect 1409 1102 1478 1107
rect 1505 1102 1550 1107
rect 1601 1102 1638 1107
rect 1777 1102 1926 1107
rect 1265 1097 1390 1102
rect 1657 1097 1758 1102
rect 297 1092 414 1097
rect 489 1092 518 1097
rect 545 1092 926 1097
rect 953 1092 1270 1097
rect 1385 1092 1430 1097
rect 1441 1092 1662 1097
rect 1753 1092 1902 1097
rect 409 1087 494 1092
rect 1425 1087 1430 1092
rect 585 1082 702 1087
rect 833 1082 966 1087
rect 1097 1082 1390 1087
rect 1425 1082 1534 1087
rect 1553 1082 1942 1087
rect 985 1077 1078 1082
rect 73 1072 174 1077
rect 489 1072 742 1077
rect 809 1072 990 1077
rect 1073 1072 1510 1077
rect 1521 1072 1790 1077
rect 385 1062 494 1067
rect 489 1057 494 1062
rect 569 1062 598 1067
rect 641 1062 910 1067
rect 945 1062 1158 1067
rect 1177 1062 1798 1067
rect 569 1057 574 1062
rect 945 1057 950 1062
rect 0 1052 102 1057
rect 201 1052 302 1057
rect 337 1052 422 1057
rect 489 1052 574 1057
rect 705 1052 950 1057
rect 961 1052 1214 1057
rect 1241 1052 1526 1057
rect 1537 1052 1590 1057
rect 1609 1052 1726 1057
rect 1809 1052 1934 1057
rect 97 1037 102 1052
rect 345 1042 374 1047
rect 393 1042 470 1047
rect 721 1042 758 1047
rect 769 1042 830 1047
rect 961 1042 966 1052
rect 1721 1047 1814 1052
rect 1001 1042 1030 1047
rect 1041 1042 1102 1047
rect 1145 1042 1702 1047
rect 849 1037 966 1042
rect 0 1032 78 1037
rect 97 1032 174 1037
rect 217 1032 278 1037
rect 353 1032 438 1037
rect 545 1032 598 1037
rect 697 1032 854 1037
rect 977 1032 1062 1037
rect 1153 1032 1222 1037
rect 1257 1032 1774 1037
rect 169 1027 174 1032
rect 1217 1027 1222 1032
rect 169 1022 342 1027
rect 449 1022 534 1027
rect 617 1022 646 1027
rect 769 1022 838 1027
rect 873 1022 894 1027
rect 945 1022 1046 1027
rect 1073 1022 1142 1027
rect 1161 1022 1206 1027
rect 1217 1022 1254 1027
rect 337 1017 454 1022
rect 529 1017 622 1022
rect 1201 1017 1206 1022
rect 113 1012 158 1017
rect 257 1012 294 1017
rect 673 1012 958 1017
rect 985 1012 1030 1017
rect 1049 1012 1110 1017
rect 1121 1012 1150 1017
rect 1201 1012 1238 1017
rect 297 1002 318 1007
rect 329 1002 430 1007
rect 497 1002 598 1007
rect 625 1002 686 1007
rect 697 1002 758 1007
rect 785 1002 974 1007
rect 985 1002 1134 1007
rect 1185 1002 1254 1007
rect 129 992 190 997
rect 225 992 286 997
rect 321 992 374 997
rect 385 992 494 997
rect 553 992 622 997
rect 641 992 678 997
rect 697 992 1262 997
rect 73 982 102 987
rect 185 982 318 987
rect 337 982 398 987
rect 433 982 478 987
rect 657 982 790 987
rect 801 982 918 987
rect 953 982 1014 987
rect 1049 982 1126 987
rect 1201 982 1270 987
rect 1281 982 1286 1027
rect 1385 1022 1558 1027
rect 1577 1022 1638 1027
rect 1649 1022 1686 1027
rect 1705 1022 1798 1027
rect 1913 1022 1950 1027
rect 1649 1017 1654 1022
rect 1793 1017 1798 1022
rect 1297 997 1302 1017
rect 1377 1012 1398 1017
rect 1457 1012 1486 1017
rect 1521 1012 1574 1017
rect 1585 1012 1654 1017
rect 1697 1012 1758 1017
rect 1793 1012 1838 1017
rect 1377 1002 1382 1012
rect 1457 1007 1462 1012
rect 1457 1002 1502 1007
rect 1297 992 1318 997
rect 1329 992 1446 997
rect 1513 992 1638 997
rect 1649 992 1686 997
rect 1329 987 1334 992
rect 1441 987 1518 992
rect 1649 987 1654 992
rect 1697 987 1702 1012
rect 1857 1007 1862 1017
rect 1857 1002 1894 1007
rect 1737 992 1758 997
rect 1769 992 1934 997
rect 1297 982 1334 987
rect 1361 982 1382 987
rect 1609 982 1654 987
rect 1673 982 1702 987
rect 1841 982 1918 987
rect 97 977 190 982
rect 265 972 422 977
rect 433 967 438 982
rect 473 977 662 982
rect 1721 977 1846 982
rect 681 972 1374 977
rect 1505 972 1726 977
rect 1857 972 1910 977
rect 137 962 230 967
rect 313 962 438 967
rect 553 962 646 967
rect 553 957 558 962
rect 0 952 78 957
rect 153 952 406 957
rect 417 952 446 957
rect 529 952 558 957
rect 641 957 646 962
rect 689 962 798 967
rect 817 962 878 967
rect 953 962 1006 967
rect 1065 962 1262 967
rect 1281 962 1334 967
rect 1393 962 1462 967
rect 1617 962 2014 967
rect 689 957 694 962
rect 641 952 694 957
rect 769 952 950 957
rect 964 952 1022 957
rect 1049 952 1238 957
rect 1321 952 1358 957
rect 1385 952 1470 957
rect 1505 952 1630 957
rect 1681 952 1782 957
rect 1801 952 1830 957
rect 1873 952 1902 957
rect 1913 952 1958 957
rect 121 942 174 947
rect 193 942 238 947
rect 273 942 334 947
rect 569 942 638 947
rect 657 942 782 947
rect 817 942 870 947
rect 905 942 934 947
rect 129 932 246 937
rect 281 932 318 937
rect 401 932 470 937
rect 513 932 614 937
rect 249 922 294 927
rect 377 922 494 927
rect 617 922 638 927
rect 153 917 230 922
rect 657 917 662 942
rect 689 932 734 937
rect 761 932 814 937
rect 897 932 942 937
rect 777 922 806 927
rect 801 917 806 922
rect 913 922 958 927
rect 913 917 918 922
rect 964 917 969 952
rect 1233 947 1326 952
rect 1113 942 1214 947
rect 1345 942 1454 947
rect 1161 932 1246 937
rect 1489 927 1494 947
rect 1521 942 1598 947
rect 1649 942 1686 947
rect 1665 932 1694 937
rect 1665 927 1670 932
rect 977 922 1054 927
rect 1081 922 1174 927
rect 1209 922 1302 927
rect 1345 922 1422 927
rect 1465 922 1494 927
rect 1521 922 1558 927
rect 1569 922 1630 927
rect 1649 922 1670 927
rect 1777 922 1782 952
rect 1825 947 1830 952
rect 1793 922 1798 947
rect 1825 942 1886 947
rect 1873 932 1894 937
rect 1889 922 1894 932
rect 1937 927 1942 947
rect 1921 922 1942 927
rect 1521 917 1526 922
rect 73 912 158 917
rect 225 912 366 917
rect 401 912 446 917
rect 609 912 662 917
rect 681 912 750 917
rect 801 912 918 917
rect 937 912 969 917
rect 977 912 1526 917
rect 1553 912 1774 917
rect 1865 912 1918 917
rect 609 907 614 912
rect 1953 907 1958 952
rect 169 902 198 907
rect 217 902 350 907
rect 417 902 614 907
rect 625 902 654 907
rect 953 902 1046 907
rect 1121 902 1238 907
rect 1281 902 1326 907
rect 1345 902 1366 907
rect 1377 902 1502 907
rect 1593 902 1662 907
rect 1673 902 1718 907
rect 1905 902 1958 907
rect 1361 897 1366 902
rect 185 892 270 897
rect 281 892 318 897
rect 945 892 1150 897
rect 1161 892 1342 897
rect 1361 892 1582 897
rect 1601 892 1790 897
rect 137 882 238 887
rect 369 882 438 887
rect 1009 882 1230 887
rect 1313 882 1398 887
rect 1393 877 1398 882
rect 1497 882 1542 887
rect 1585 882 1838 887
rect 1497 877 1502 882
rect 0 872 78 877
rect 929 872 1294 877
rect 1393 872 1502 877
rect 1537 872 1662 877
rect 1697 872 1758 877
rect 1769 872 1910 877
rect 1697 867 1702 872
rect 305 862 374 867
rect 305 857 310 862
rect 0 852 310 857
rect 369 857 374 862
rect 529 862 614 867
rect 1001 862 1110 867
rect 1241 862 1374 867
rect 1521 862 1702 867
rect 1713 862 1854 867
rect 529 857 534 862
rect 369 852 398 857
rect 505 852 534 857
rect 609 857 614 862
rect 1129 857 1222 862
rect 609 852 710 857
rect 937 852 1134 857
rect 1217 852 1478 857
rect 1529 852 1566 857
rect 1697 852 1750 857
rect 1585 847 1702 852
rect 321 842 462 847
rect 777 842 910 847
rect 929 842 1278 847
rect 1305 842 1366 847
rect 1441 842 1590 847
rect 1721 842 1878 847
rect 777 837 782 842
rect 225 832 254 837
rect 377 832 422 837
rect 433 832 598 837
rect 721 832 782 837
rect 905 837 910 842
rect 905 832 942 837
rect 985 832 1030 837
rect 1041 832 1126 837
rect 1145 832 1166 837
rect 1177 832 1214 837
rect 1281 832 1438 837
rect 1473 832 1774 837
rect 1801 832 1862 837
rect 433 827 438 832
rect 193 822 302 827
rect 329 822 438 827
rect 449 822 494 827
rect 569 822 678 827
rect 873 822 902 827
rect 945 822 998 827
rect 73 812 358 817
rect 409 812 518 817
rect 585 812 638 817
rect 665 812 710 817
rect 793 812 862 817
rect 889 812 950 817
rect 513 807 518 812
rect 177 802 198 807
rect 273 802 342 807
rect 361 802 438 807
rect 513 802 566 807
rect 593 802 958 807
rect 297 792 326 797
rect 561 792 614 797
rect 625 792 670 797
rect 681 792 726 797
rect 769 792 830 797
rect 841 792 878 797
rect 897 792 966 797
rect 409 787 534 792
rect 993 787 998 822
rect 1025 807 1030 832
rect 1089 822 1126 827
rect 1137 822 1246 827
rect 1273 822 1318 827
rect 1121 817 1126 822
rect 1057 812 1102 817
rect 1121 812 1334 817
rect 1025 802 1062 807
rect 1081 802 1294 807
rect 1393 797 1398 827
rect 1417 822 1446 827
rect 1457 822 1633 827
rect 1441 807 1446 822
rect 1628 817 1633 822
rect 1641 817 1646 827
rect 1689 822 1742 827
rect 1441 802 1478 807
rect 1073 792 1398 797
rect 225 782 254 787
rect 385 782 414 787
rect 529 782 558 787
rect 705 782 982 787
rect 993 782 1030 787
rect 1105 782 1286 787
rect 1305 782 1374 787
rect 1385 782 1422 787
rect 1441 782 1494 787
rect 1105 777 1110 782
rect 1505 777 1510 817
rect 1521 802 1598 807
rect 1521 782 1526 802
rect 1617 797 1622 817
rect 1628 812 1638 817
rect 1641 812 1654 817
rect 1713 812 1742 817
rect 1593 792 1622 797
rect 1633 787 1638 812
rect 1649 807 1654 812
rect 1649 802 1670 807
rect 1657 792 1750 797
rect 1537 782 1574 787
rect 1633 782 1710 787
rect 209 772 278 777
rect 425 772 518 777
rect 553 772 694 777
rect 753 772 830 777
rect 969 772 1110 777
rect 1121 772 1150 777
rect 1217 772 1302 777
rect 1313 772 1646 777
rect 689 767 694 772
rect 1297 767 1302 772
rect 265 762 438 767
rect 521 762 550 767
rect 617 762 670 767
rect 689 762 718 767
rect 729 762 1022 767
rect 1057 762 1142 767
rect 1169 762 1214 767
rect 1297 762 1350 767
rect 1393 762 1478 767
rect 1489 762 1678 767
rect 1697 762 1742 767
rect 0 752 70 757
rect 585 752 878 757
rect 993 752 1166 757
rect 1265 752 1334 757
rect 1345 752 1398 757
rect 145 742 174 747
rect 265 742 310 747
rect 337 742 542 747
rect 601 742 742 747
rect 753 742 814 747
rect 865 742 990 747
rect 1089 742 1150 747
rect 1161 742 1222 747
rect 225 732 254 737
rect 313 732 406 737
rect 657 732 734 737
rect 1089 727 1094 742
rect 1329 737 1334 752
rect 1153 727 1158 737
rect 129 722 198 727
rect 217 722 286 727
rect 305 722 374 727
rect 713 722 750 727
rect 769 722 790 727
rect 809 722 894 727
rect 977 722 1014 727
rect 1049 722 1094 727
rect 1105 722 1158 727
rect 1169 727 1174 737
rect 1241 732 1294 737
rect 1305 732 1334 737
rect 1361 727 1366 747
rect 1169 722 1238 727
rect 1313 722 1342 727
rect 1361 722 1382 727
rect 137 712 174 717
rect 305 707 310 722
rect 809 717 814 722
rect 377 712 430 717
rect 449 712 582 717
rect 641 712 742 717
rect 761 712 814 717
rect 889 717 894 722
rect 1009 717 1014 722
rect 1393 717 1398 752
rect 1425 727 1430 757
rect 1481 752 1518 757
rect 1537 752 1670 757
rect 1697 747 1702 762
rect 1449 742 1526 747
rect 1553 742 1622 747
rect 1633 742 1702 747
rect 1633 737 1638 742
rect 1473 732 1510 737
rect 1577 732 1638 737
rect 1425 722 1454 727
rect 1473 722 1478 732
rect 1529 722 1566 727
rect 1585 722 1630 727
rect 1641 722 1686 727
rect 1585 717 1590 722
rect 889 712 918 717
rect 945 712 998 717
rect 1009 712 1062 717
rect 1129 712 1198 717
rect 1273 712 1310 717
rect 1329 712 1374 717
rect 1393 712 1446 717
rect 1505 712 1590 717
rect 1697 717 1702 737
rect 1745 727 1750 757
rect 1729 722 1750 727
rect 1761 717 1766 827
rect 1793 822 1822 827
rect 1905 822 1990 827
rect 1777 812 1854 817
rect 1777 792 1814 797
rect 1825 792 1862 797
rect 1905 787 1910 822
rect 1921 812 1958 817
rect 1777 782 1846 787
rect 1905 782 1934 787
rect 1777 772 1854 777
rect 1865 772 1894 777
rect 1905 772 1942 777
rect 1777 727 1782 772
rect 1953 767 1958 812
rect 1985 787 1990 822
rect 1985 782 2020 787
rect 1793 762 1878 767
rect 1953 762 2020 767
rect 1793 747 1798 757
rect 1809 752 1894 757
rect 1793 742 1814 747
rect 1857 742 1926 747
rect 1777 722 1798 727
rect 1809 722 1814 742
rect 1849 732 1886 737
rect 1999 727 2004 762
rect 1999 722 2014 727
rect 1697 712 1742 717
rect 1761 712 1790 717
rect 1825 712 1862 717
rect 1873 712 2020 717
rect 449 707 454 712
rect 281 702 310 707
rect 353 702 454 707
rect 697 702 790 707
rect 825 702 1262 707
rect 1513 702 1662 707
rect 1729 702 1782 707
rect 361 692 398 697
rect 441 692 598 697
rect 785 692 1054 697
rect 1073 692 1326 697
rect 1345 692 1494 697
rect 1569 692 1670 697
rect 1705 692 1838 697
rect 1913 692 2020 697
rect 0 682 70 687
rect 217 682 342 687
rect 521 682 774 687
rect 921 682 958 687
rect 1009 682 1014 692
rect 1345 687 1350 692
rect 1065 682 1350 687
rect 1489 687 1494 692
rect 1489 682 1758 687
rect 769 677 902 682
rect 1817 677 1918 682
rect 105 672 350 677
rect 425 672 566 677
rect 897 672 1230 677
rect 585 667 734 672
rect 1225 667 1230 672
rect 1329 672 1694 677
rect 1793 672 1822 677
rect 1913 672 2020 677
rect 1329 667 1334 672
rect 265 662 318 667
rect 361 662 454 667
rect 561 662 590 667
rect 729 662 758 667
rect 769 662 942 667
rect 1025 662 1078 667
rect 1137 662 1206 667
rect 1225 662 1334 667
rect 1441 662 1518 667
rect 1729 662 1934 667
rect 1537 657 1710 662
rect 169 652 534 657
rect 585 652 1070 657
rect 1081 652 1190 657
rect 1401 652 1542 657
rect 1705 652 1846 657
rect 185 642 214 647
rect 289 642 334 647
rect 609 642 646 647
rect 729 642 878 647
rect 897 642 974 647
rect 985 642 1030 647
rect 1153 642 1270 647
rect 1337 642 1766 647
rect 1777 642 1934 647
rect 441 637 590 642
rect 137 632 446 637
rect 585 632 774 637
rect 881 632 902 637
rect 929 632 1006 637
rect 1129 632 1206 637
rect 1217 632 1318 637
rect 1329 632 1486 637
rect 1545 632 1582 637
rect 1201 627 1206 632
rect 1329 627 1334 632
rect 1681 627 1774 632
rect 65 617 70 627
rect 113 622 206 627
rect 257 622 278 627
rect 321 622 390 627
rect 457 622 606 627
rect 65 612 86 617
rect 81 607 86 612
rect 185 612 222 617
rect 185 607 190 612
rect 81 602 190 607
rect 273 607 278 622
rect 297 612 382 617
rect 521 612 558 617
rect 593 612 638 617
rect 273 602 302 607
rect 329 602 398 607
rect 569 602 614 607
rect 625 602 734 607
rect 241 592 270 597
rect 313 592 342 597
rect 337 587 342 592
rect 409 592 446 597
rect 513 592 582 597
rect 617 592 678 597
rect 409 587 414 592
rect 209 582 318 587
rect 337 582 414 587
rect 465 582 566 587
rect 577 582 646 587
rect 753 582 758 627
rect 841 622 894 627
rect 977 622 1062 627
rect 1097 622 1142 627
rect 1201 622 1334 627
rect 1345 622 1430 627
rect 1465 622 1510 627
rect 1553 622 1606 627
rect 1657 622 1686 627
rect 1769 622 1798 627
rect 1817 622 1870 627
rect 1881 622 1918 627
rect 1793 617 1798 622
rect 769 577 774 617
rect 873 612 1358 617
rect 1377 612 1406 617
rect 1497 612 1526 617
rect 1377 607 1382 612
rect 841 602 1022 607
rect 1193 602 1270 607
rect 1361 602 1382 607
rect 1449 602 1478 607
rect 1041 597 1174 602
rect 905 592 966 597
rect 985 592 1046 597
rect 1169 592 1342 597
rect 1353 592 1502 597
rect 1521 592 1526 612
rect 1537 607 1542 617
rect 1585 612 1718 617
rect 1537 602 1566 607
rect 1665 602 1702 607
rect 1561 597 1670 602
rect 1713 597 1718 612
rect 1689 592 1718 597
rect 1729 587 1734 617
rect 1753 612 1782 617
rect 1793 612 1950 617
rect 1777 597 1782 612
rect 1969 602 2020 607
rect 1761 592 1782 597
rect 1833 592 1934 597
rect 1969 587 1974 602
rect 953 582 1134 587
rect 1145 582 1190 587
rect 1201 582 1318 587
rect 1401 582 1462 587
rect 1489 582 1734 587
rect 1769 582 1974 587
rect 217 572 294 577
rect 545 572 654 577
rect 745 572 806 577
rect 881 572 990 577
rect 1001 572 1126 577
rect 1153 572 1246 577
rect 1329 572 1614 577
rect 1657 572 1886 577
rect 1929 572 2020 577
rect 1153 567 1158 572
rect 1241 567 1334 572
rect 129 562 190 567
rect 273 562 310 567
rect 473 562 894 567
rect 977 562 1158 567
rect 1169 562 1222 567
rect 1369 562 1486 567
rect 1625 562 1878 567
rect 1481 557 1630 562
rect 233 552 326 557
rect 409 552 454 557
rect 481 552 502 557
rect 625 552 678 557
rect 137 542 246 547
rect 255 542 270 547
rect 441 542 470 547
rect 255 537 260 542
rect 121 532 174 537
rect 225 532 260 537
rect 273 532 334 537
rect 105 512 206 517
rect 73 502 214 507
rect 225 502 230 532
rect 481 527 486 552
rect 529 542 638 547
rect 649 542 678 547
rect 329 522 454 527
rect 465 522 486 527
rect 497 532 558 537
rect 641 532 662 537
rect 497 522 502 532
rect 561 522 630 527
rect 641 522 646 532
rect 673 522 678 542
rect 689 527 694 557
rect 721 552 750 557
rect 785 547 790 557
rect 913 552 1094 557
rect 1185 552 1214 557
rect 721 542 790 547
rect 841 542 910 547
rect 929 542 958 547
rect 969 542 1206 547
rect 929 537 934 542
rect 729 532 934 537
rect 977 532 1046 537
rect 1113 532 1182 537
rect 1041 527 1046 532
rect 1233 527 1238 557
rect 1257 552 1366 557
rect 1441 552 1462 557
rect 1665 552 1822 557
rect 1833 552 1862 557
rect 1249 542 1350 547
rect 1377 542 1430 547
rect 1329 532 1358 537
rect 1441 527 1446 552
rect 1665 547 1670 552
rect 1833 547 1838 552
rect 1481 542 1582 547
rect 1601 542 1670 547
rect 1681 542 1750 547
rect 1761 542 1838 547
rect 1481 537 1486 542
rect 689 522 910 527
rect 1041 522 1118 527
rect 1217 522 1238 527
rect 1401 522 1446 527
rect 1457 532 1486 537
rect 1577 537 1582 542
rect 1857 537 1862 552
rect 1897 552 1974 557
rect 1897 547 1902 552
rect 1873 542 1902 547
rect 1969 547 1974 552
rect 1969 542 2014 547
rect 1577 532 1830 537
rect 1857 532 1958 537
rect 249 512 318 517
rect 345 512 390 517
rect 401 512 446 517
rect 481 512 598 517
rect 617 512 662 517
rect 681 512 886 517
rect 897 512 966 517
rect 977 512 1030 517
rect 1081 512 1110 517
rect 1137 512 1238 517
rect 1257 512 1294 517
rect 1305 512 1382 517
rect 1393 512 1430 517
rect 401 507 406 512
rect 593 507 598 512
rect 1377 507 1382 512
rect 1457 507 1462 532
rect 1513 522 1630 527
rect 1761 522 1798 527
rect 1809 522 1846 527
rect 1625 517 1766 522
rect 1545 512 1598 517
rect 1785 512 1830 517
rect 1841 507 1846 522
rect 1953 517 1958 532
rect 1913 512 1958 517
rect 241 502 262 507
rect 289 502 406 507
rect 449 502 502 507
rect 513 502 566 507
rect 593 502 830 507
rect 849 502 990 507
rect 1033 502 1078 507
rect 1097 502 1270 507
rect 1281 502 1318 507
rect 1377 502 1462 507
rect 1505 502 1574 507
rect 1649 502 1822 507
rect 1841 502 1934 507
rect 241 497 246 502
rect 513 497 518 502
rect 1265 497 1270 502
rect 169 492 246 497
rect 265 492 398 497
rect 441 492 518 497
rect 593 492 918 497
rect 969 492 1142 497
rect 1161 492 1238 497
rect 1265 492 1422 497
rect 1433 492 1494 497
rect 1513 492 1582 497
rect 1753 492 1854 497
rect 1233 487 1238 492
rect 1849 487 1854 492
rect 1969 492 2014 497
rect 1969 487 1974 492
rect 0 482 262 487
rect 337 482 1222 487
rect 1233 482 1310 487
rect 1321 482 1462 487
rect 1561 482 1694 487
rect 1721 482 1758 487
rect 1849 482 1974 487
rect 113 472 222 477
rect 433 472 1030 477
rect 1041 472 1150 477
rect 1185 472 1526 477
rect 1681 472 1830 477
rect 1041 467 1046 472
rect 81 462 334 467
rect 465 462 550 467
rect 561 462 646 467
rect 673 462 1046 467
rect 1057 462 1142 467
rect 1153 462 1782 467
rect 353 457 446 462
rect 153 452 198 457
rect 321 452 358 457
rect 441 452 774 457
rect 881 452 1094 457
rect 1105 452 1182 457
rect 1193 452 1438 457
rect 1649 452 1886 457
rect 769 447 886 452
rect 1433 447 1558 452
rect 1649 447 1654 452
rect 377 442 446 447
rect 473 442 526 447
rect 545 442 614 447
rect 625 442 750 447
rect 905 442 1158 447
rect 1169 442 1214 447
rect 1225 442 1326 447
rect 1345 442 1414 447
rect 1553 442 1654 447
rect 1705 442 1814 447
rect 289 432 414 437
rect 473 432 510 437
rect 553 432 590 437
rect 153 422 230 427
rect 313 422 358 427
rect 401 422 446 427
rect 489 422 550 427
rect 561 422 606 427
rect 225 417 230 422
rect 545 417 550 422
rect 97 412 182 417
rect 225 412 366 417
rect 417 412 438 417
rect 449 412 470 417
rect 97 387 102 412
rect 433 407 438 412
rect 353 402 382 407
rect 409 402 438 407
rect 465 402 470 412
rect 529 407 534 417
rect 545 412 574 417
rect 625 407 630 442
rect 1809 437 1814 442
rect 1889 442 1918 447
rect 1889 437 1894 442
rect 529 402 566 407
rect 577 402 630 407
rect 641 432 710 437
rect 721 432 814 437
rect 833 432 902 437
rect 913 432 1030 437
rect 1057 432 1102 437
rect 1113 432 1406 437
rect 1417 432 1534 437
rect 1673 432 1702 437
rect 177 392 198 397
rect 257 392 310 397
rect 417 392 502 397
rect 545 392 598 397
rect 0 382 102 387
rect 209 382 334 387
rect 393 382 510 387
rect 641 382 646 432
rect 833 427 838 432
rect 897 427 902 432
rect 721 422 774 427
rect 801 422 838 427
rect 849 422 886 427
rect 897 422 966 427
rect 993 422 1022 427
rect 657 412 686 417
rect 721 412 726 422
rect 1057 417 1062 432
rect 1081 422 1142 427
rect 657 392 662 412
rect 737 407 742 417
rect 785 407 790 417
rect 897 412 942 417
rect 953 412 1062 417
rect 1097 412 1134 417
rect 673 402 742 407
rect 753 402 790 407
rect 993 402 1118 407
rect 673 387 678 402
rect 809 397 950 402
rect 1153 397 1158 427
rect 1185 402 1190 432
rect 1217 412 1238 417
rect 1233 402 1238 412
rect 1249 397 1254 427
rect 705 392 750 397
rect 769 392 814 397
rect 945 392 1006 397
rect 1065 392 1102 397
rect 1153 392 1198 397
rect 1217 392 1254 397
rect 1265 397 1270 427
rect 1281 422 1374 427
rect 1385 422 1406 427
rect 1433 422 1510 427
rect 1601 422 1694 427
rect 1297 397 1302 417
rect 1481 407 1574 412
rect 1321 402 1414 407
rect 1457 402 1486 407
rect 1569 402 1598 407
rect 1321 397 1326 402
rect 1265 392 1286 397
rect 1297 392 1326 397
rect 1409 397 1414 402
rect 1649 397 1654 417
rect 1665 412 1686 417
rect 1409 392 1438 397
rect 1481 392 1670 397
rect 769 387 774 392
rect 657 382 678 387
rect 689 382 718 387
rect 737 382 774 387
rect 817 382 958 387
rect 1009 382 1582 387
rect 241 372 326 377
rect 537 372 782 377
rect 857 372 998 377
rect 121 367 222 372
rect 1009 367 1014 382
rect 1681 377 1686 412
rect 1729 387 1734 417
rect 1745 407 1750 437
rect 1761 432 1790 437
rect 1809 432 1894 437
rect 1745 402 1766 407
rect 1713 382 1734 387
rect 1777 382 1782 427
rect 1793 412 1814 417
rect 1809 392 1814 412
rect 1889 407 1894 417
rect 1833 402 1918 407
rect 1841 392 1942 397
rect 1849 382 1894 387
rect 1057 372 1078 377
rect 1105 372 1166 377
rect 1177 372 1206 377
rect 1265 372 1534 377
rect 1633 372 1662 377
rect 1681 372 1766 377
rect 0 362 126 367
rect 217 362 310 367
rect 401 362 430 367
rect 489 362 558 367
rect 585 362 654 367
rect 697 362 734 367
rect 753 362 798 367
rect 961 362 1014 367
rect 1033 362 1078 367
rect 1121 362 1254 367
rect 1273 362 1406 367
rect 1433 362 1502 367
rect 1721 362 1950 367
rect 961 357 966 362
rect 137 352 254 357
rect 561 352 966 357
rect 145 342 270 347
rect 289 342 374 347
rect 417 342 462 347
rect 481 342 526 347
rect 609 342 694 347
rect 713 342 774 347
rect 833 342 862 347
rect 609 337 614 342
rect 465 332 614 337
rect 689 337 694 342
rect 689 332 790 337
rect 841 327 942 332
rect 201 322 238 327
rect 265 322 302 327
rect 401 322 430 327
rect 449 322 494 327
rect 601 322 646 327
rect 665 322 710 327
rect 737 322 798 327
rect 817 322 846 327
rect 937 322 966 327
rect 977 322 982 357
rect 1001 347 1006 357
rect 1025 352 1062 357
rect 993 342 1006 347
rect 993 327 998 342
rect 1057 337 1062 352
rect 1073 347 1078 362
rect 1089 352 1142 357
rect 1153 352 1190 357
rect 1377 352 1446 357
rect 1465 352 1510 357
rect 1641 352 1702 357
rect 1745 352 1814 357
rect 1073 342 1126 347
rect 1153 342 1214 347
rect 1225 342 1262 347
rect 1281 342 1638 347
rect 1649 342 1782 347
rect 1809 342 1838 347
rect 1281 337 1286 342
rect 1057 332 1078 337
rect 1073 327 1078 332
rect 1161 332 1286 337
rect 1337 332 1374 337
rect 1409 332 1454 337
rect 1161 327 1166 332
rect 993 322 1054 327
rect 1073 322 1166 327
rect 1473 327 1478 337
rect 1633 327 1638 342
rect 1657 332 1694 337
rect 1473 322 1558 327
rect 1633 322 1750 327
rect 1809 322 1814 342
rect 1857 322 1894 327
rect 737 317 742 322
rect 961 317 966 322
rect 1209 317 1278 322
rect 1345 317 1422 322
rect 1857 317 1862 322
rect 249 312 318 317
rect 353 312 590 317
rect 697 312 742 317
rect 777 312 886 317
rect 905 312 942 317
rect 961 312 1046 317
rect 1185 312 1214 317
rect 1273 312 1350 317
rect 1417 312 1446 317
rect 1473 312 1534 317
rect 1673 312 1742 317
rect 1833 312 1862 317
rect 1441 307 1446 312
rect 1905 307 1910 357
rect 217 302 294 307
rect 369 302 422 307
rect 457 302 502 307
rect 513 302 822 307
rect 873 302 934 307
rect 945 302 982 307
rect 1137 302 1262 307
rect 1361 302 1422 307
rect 1441 302 1470 307
rect 1545 302 1662 307
rect 1737 302 1862 307
rect 1881 302 1910 307
rect 1465 297 1550 302
rect 1657 297 1742 302
rect 257 292 334 297
rect 441 292 534 297
rect 585 292 830 297
rect 889 292 942 297
rect 1217 292 1270 297
rect 1761 292 1846 297
rect 329 282 390 287
rect 457 282 846 287
rect 857 282 918 287
rect 1001 282 1118 287
rect 1457 282 1750 287
rect 1857 282 1942 287
rect 1001 277 1006 282
rect 353 272 894 277
rect 905 272 1006 277
rect 1113 277 1118 282
rect 1745 277 1862 282
rect 1113 272 1190 277
rect 1233 272 1286 277
rect 1297 272 1486 277
rect 1481 267 1486 272
rect 1593 272 1622 277
rect 1593 267 1598 272
rect 393 262 462 267
rect 577 262 782 267
rect 897 262 1142 267
rect 1201 262 1278 267
rect 1481 262 1598 267
rect 1745 262 1862 267
rect 433 252 478 257
rect 601 252 622 257
rect 633 252 670 257
rect 841 252 974 257
rect 1193 252 1350 257
rect 1817 252 1918 257
rect 1105 247 1174 252
rect 313 242 790 247
rect 801 242 1110 247
rect 1169 242 1462 247
rect 1673 242 1814 247
rect 801 237 806 242
rect 73 232 230 237
rect 473 232 806 237
rect 825 232 950 237
rect 1121 232 1334 237
rect 1449 232 1486 237
rect 1705 232 1742 237
rect 289 222 382 227
rect 401 222 446 227
rect 465 222 542 227
rect 561 222 614 227
rect 665 222 766 227
rect 817 222 854 227
rect 865 222 902 227
rect 929 222 1006 227
rect 1017 222 1102 227
rect 1137 222 1166 227
rect 1233 222 1278 227
rect 1337 222 1366 227
rect 1377 222 1422 227
rect 1441 222 1558 227
rect 1609 222 1638 227
rect 1721 222 1750 227
rect 401 217 406 222
rect 193 212 230 217
rect 273 212 310 217
rect 361 212 406 217
rect 465 207 470 222
rect 489 212 558 217
rect 585 212 646 217
rect 673 212 742 217
rect 777 212 894 217
rect 921 212 1014 217
rect 1049 212 1110 217
rect 313 202 470 207
rect 529 202 638 207
rect 689 202 734 207
rect 785 202 830 207
rect 849 202 886 207
rect 1057 202 1094 207
rect 153 192 198 197
rect 225 192 502 197
rect 673 192 798 197
rect 849 192 854 202
rect 1105 197 1110 212
rect 1137 207 1142 222
rect 1377 217 1382 222
rect 1153 212 1310 217
rect 1329 212 1382 217
rect 1425 212 1542 217
rect 1633 207 1638 222
rect 1657 212 1702 217
rect 1137 202 1182 207
rect 1257 202 1318 207
rect 1633 202 1678 207
rect 1001 192 1078 197
rect 1105 192 1126 197
rect 1289 192 1326 197
rect 1337 192 1454 197
rect 1473 192 1542 197
rect 1593 192 1734 197
rect 1473 187 1478 192
rect 217 182 286 187
rect 321 182 414 187
rect 457 182 486 187
rect 505 182 590 187
rect 617 182 678 187
rect 721 182 878 187
rect 889 182 974 187
rect 985 182 1206 187
rect 1281 182 1478 187
rect 1537 187 1542 192
rect 1537 182 1670 187
rect 1745 182 1750 222
rect 1793 217 1798 227
rect 1761 212 1798 217
rect 1809 197 1814 242
rect 1873 222 1918 227
rect 1793 192 1814 197
rect 1857 192 1862 217
rect 1897 212 1934 217
rect 1793 177 1798 192
rect 1809 182 1846 187
rect 465 172 582 177
rect 753 167 758 177
rect 801 172 1246 177
rect 1265 172 1318 177
rect 1329 172 1382 177
rect 1433 172 1462 177
rect 1473 172 1526 177
rect 1705 172 1734 177
rect 1777 172 1798 177
rect 1817 172 1854 177
rect 1777 167 1782 172
rect 385 162 438 167
rect 449 162 526 167
rect 601 162 702 167
rect 737 162 830 167
rect 857 162 886 167
rect 1073 162 1174 167
rect 1209 162 1246 167
rect 1297 162 1430 167
rect 1601 162 1654 167
rect 1705 162 1782 167
rect 1793 162 1830 167
rect 1849 162 1878 167
rect 601 157 606 162
rect 289 152 334 157
rect 345 152 606 157
rect 697 157 702 162
rect 905 157 1054 162
rect 697 152 726 157
rect 857 152 910 157
rect 1049 152 1094 157
rect 1177 152 1294 157
rect 1465 152 1550 157
rect 721 147 862 152
rect 1089 147 1182 152
rect 1313 147 1446 152
rect 1745 147 1750 157
rect 1833 152 1886 157
rect 369 142 430 147
rect 497 142 566 147
rect 609 142 686 147
rect 561 137 566 142
rect 881 137 886 147
rect 945 142 982 147
rect 1033 142 1070 147
rect 1201 142 1318 147
rect 1441 142 1502 147
rect 1561 142 1782 147
rect 1793 142 1862 147
rect 1497 137 1566 142
rect 561 132 606 137
rect 625 132 766 137
rect 817 127 822 137
rect 417 122 510 127
rect 793 122 822 127
rect 849 132 886 137
rect 257 112 278 117
rect 289 112 342 117
rect 529 112 630 117
rect 769 112 822 117
rect 849 112 854 132
rect 1121 127 1126 137
rect 1185 127 1190 137
rect 1217 132 1302 137
rect 1313 132 1478 137
rect 1473 127 1478 132
rect 1121 122 1150 127
rect 1185 122 1214 127
rect 1377 122 1414 127
rect 1425 122 1462 127
rect 1473 122 1582 127
rect 1657 122 1726 127
rect 1913 122 1934 127
rect 977 112 1062 117
rect 1177 112 1222 117
rect 1281 112 1350 117
rect 1401 112 1446 117
rect 1457 112 1462 122
rect 1553 112 1646 117
rect 1665 112 1894 117
rect 305 102 414 107
rect 425 102 518 107
rect 617 102 758 107
rect 857 102 910 107
rect 1129 102 1190 107
rect 1249 102 1406 107
rect 1417 102 1534 107
rect 1609 102 1686 107
rect 753 97 862 102
rect 425 92 550 97
rect 881 92 1198 97
rect 1209 92 1270 97
rect 1313 92 1358 97
rect 1473 92 1638 97
rect 1353 87 1478 92
rect 497 82 958 87
rect 1201 82 1334 87
rect 1329 77 1334 82
rect 1497 82 1526 87
rect 1497 77 1502 82
rect 681 72 710 77
rect 705 67 710 72
rect 945 72 1126 77
rect 1265 72 1310 77
rect 1329 72 1502 77
rect 1649 72 1790 77
rect 945 67 950 72
rect 705 62 950 67
rect 969 62 1254 67
rect 1305 57 1310 72
rect 1649 67 1654 72
rect 1537 62 1654 67
rect 1537 57 1542 62
rect 1145 52 1286 57
rect 1305 52 1542 57
rect 1041 47 1126 52
rect 745 42 942 47
rect 961 42 1046 47
rect 1121 42 1190 47
rect 745 27 750 42
rect 593 22 750 27
rect 937 27 942 42
rect 1057 32 1222 37
rect 937 22 1206 27
rect 761 12 926 17
rect 921 7 926 12
rect 1057 12 1134 17
rect 1361 12 1398 17
rect 1057 7 1062 12
rect 921 2 1062 7
use top_module_VIA1  top_module_VIA1_0
timestamp 1524952243
transform 1 0 24 0 1 1917
box -10 -10 10 10
use M3_M2  M3_M2_0
timestamp 1524952243
transform 1 0 1300 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1524952243
transform 1 0 1324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1524952243
transform 1 0 1332 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1524952243
transform 1 0 1396 0 1 1915
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1524952243
transform 1 0 48 0 1 1893
box -10 -10 10 10
use M3_M2  M3_M2_4
timestamp 1524952243
transform 1 0 972 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1524952243
transform 1 0 1068 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1524952243
transform 1 0 1396 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1524952243
transform 1 0 1444 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1524952243
transform 1 0 1524 0 1 1905
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1524952243
transform 1 0 1994 0 1 1917
box -10 -10 10 10
use M3_M2  M3_M2_9
timestamp 1524952243
transform 1 0 956 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1524952243
transform 1 0 1052 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1524952243
transform 1 0 940 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1524952243
transform 1 0 1084 0 1 1885
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1524952243
transform 1 0 1970 0 1 1893
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_0
timestamp 1524952243
transform 1 0 24 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_36
timestamp 1524952243
transform 1 0 180 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_22
timestamp 1524952243
transform 1 0 76 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1524952243
transform 1 0 84 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1524952243
transform 1 0 132 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1524952243
transform 1 0 172 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_24
timestamp 1524952243
transform 1 0 180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1524952243
transform 1 0 156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1524952243
transform 1 0 172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1524952243
transform 1 0 132 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1524952243
transform 1 0 212 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1524952243
transform 1 0 212 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_0
timestamp 1524952243
transform 1 0 252 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1524952243
transform 1 0 244 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1524952243
transform 1 0 228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1524952243
transform 1 0 204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1524952243
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1524952243
transform 1 0 212 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1524952243
transform 1 0 268 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1524952243
transform 1 0 292 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1
timestamp 1524952243
transform 1 0 332 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1524952243
transform 1 0 308 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1524952243
transform 1 0 332 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1524952243
transform 1 0 260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1524952243
transform 1 0 276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1524952243
transform 1 0 292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1524952243
transform 1 0 300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1524952243
transform 1 0 308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1524952243
transform 1 0 236 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1524952243
transform 1 0 260 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1524952243
transform 1 0 276 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_88
timestamp 1524952243
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_121
timestamp 1524952243
transform 1 0 284 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1524952243
transform 1 0 308 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1524952243
transform 1 0 340 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1524952243
transform 1 0 356 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1524952243
transform 1 0 340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1524952243
transform 1 0 364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1524952243
transform 1 0 404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1524952243
transform 1 0 324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1524952243
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1524952243
transform 1 0 364 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1524952243
transform 1 0 404 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_34
timestamp 1524952243
transform 1 0 508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1524952243
transform 1 0 548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1524952243
transform 1 0 572 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_74
timestamp 1524952243
transform 1 0 580 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_91
timestamp 1524952243
transform 1 0 468 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1524952243
transform 1 0 508 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1524952243
transform 1 0 532 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1524952243
transform 1 0 548 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_92
timestamp 1524952243
transform 1 0 556 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_90
timestamp 1524952243
transform 1 0 580 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1524952243
transform 1 0 612 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1524952243
transform 1 0 604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1524952243
transform 1 0 612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1524952243
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1524952243
transform 1 0 652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1524952243
transform 1 0 588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1524952243
transform 1 0 596 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_106
timestamp 1524952243
transform 1 0 516 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1524952243
transform 1 0 556 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_135
timestamp 1524952243
transform 1 0 572 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1524952243
transform 1 0 604 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1524952243
transform 1 0 612 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_108
timestamp 1524952243
transform 1 0 588 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1524952243
transform 1 0 612 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_96
timestamp 1524952243
transform 1 0 644 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1524952243
transform 1 0 644 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1524952243
transform 1 0 660 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1524952243
transform 1 0 692 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1524952243
transform 1 0 676 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1524952243
transform 1 0 660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1524952243
transform 1 0 668 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_30
timestamp 1524952243
transform 1 0 732 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1524952243
transform 1 0 764 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1524952243
transform 1 0 772 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1524952243
transform 1 0 740 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1524952243
transform 1 0 756 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1524952243
transform 1 0 732 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1524952243
transform 1 0 716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1524952243
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1524952243
transform 1 0 684 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_92
timestamp 1524952243
transform 1 0 716 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1524952243
transform 1 0 756 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1524952243
transform 1 0 748 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1524952243
transform 1 0 788 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1524952243
transform 1 0 844 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1524952243
transform 1 0 828 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1524952243
transform 1 0 812 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1524952243
transform 1 0 804 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1524952243
transform 1 0 788 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1524952243
transform 1 0 772 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1524952243
transform 1 0 804 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1524952243
transform 1 0 812 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1524952243
transform 1 0 780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1524952243
transform 1 0 804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1524952243
transform 1 0 820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1524952243
transform 1 0 732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1524952243
transform 1 0 740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1524952243
transform 1 0 756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1524952243
transform 1 0 684 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_123
timestamp 1524952243
transform 1 0 684 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1524952243
transform 1 0 756 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1524952243
transform 1 0 740 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1524952243
transform 1 0 756 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_102
timestamp 1524952243
transform 1 0 780 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1524952243
transform 1 0 804 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1524952243
transform 1 0 836 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_15
timestamp 1524952243
transform 1 0 836 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_23
timestamp 1524952243
transform 1 0 868 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1524952243
transform 1 0 908 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1524952243
transform 1 0 900 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1524952243
transform 1 0 924 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1524952243
transform 1 0 892 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1524952243
transform 1 0 892 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1524952243
transform 1 0 900 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1524952243
transform 1 0 860 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1524952243
transform 1 0 876 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1524952243
transform 1 0 892 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1524952243
transform 1 0 852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1524952243
transform 1 0 836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1524952243
transform 1 0 860 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_112
timestamp 1524952243
transform 1 0 852 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_137
timestamp 1524952243
transform 1 0 868 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_31
timestamp 1524952243
transform 1 0 932 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_17
timestamp 1524952243
transform 1 0 916 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1524952243
transform 1 0 924 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1524952243
transform 1 0 884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1524952243
transform 1 0 900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1524952243
transform 1 0 884 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1524952243
transform 1 0 916 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1524952243
transform 1 0 972 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1524952243
transform 1 0 956 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_18
timestamp 1524952243
transform 1 0 940 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1524952243
transform 1 0 932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1524952243
transform 1 0 924 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1524952243
transform 1 0 964 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1524952243
transform 1 0 980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1524952243
transform 1 0 1020 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1524952243
transform 1 0 1044 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1524952243
transform 1 0 1036 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1524952243
transform 1 0 1012 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1524952243
transform 1 0 996 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1524952243
transform 1 0 956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1524952243
transform 1 0 940 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_113
timestamp 1524952243
transform 1 0 940 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1524952243
transform 1 0 1028 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1524952243
transform 1 0 980 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1524952243
transform 1 0 1004 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_54
timestamp 1524952243
transform 1 0 1028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1524952243
transform 1 0 1036 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1524952243
transform 1 0 1076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1524952243
transform 1 0 964 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1524952243
transform 1 0 972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1524952243
transform 1 0 980 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_110
timestamp 1524952243
transform 1 0 996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1524952243
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_126
timestamp 1524952243
transform 1 0 988 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1524952243
transform 1 0 1004 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1524952243
transform 1 0 1068 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_112
timestamp 1524952243
transform 1 0 1116 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_114
timestamp 1524952243
transform 1 0 1116 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1524952243
transform 1 0 1220 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1524952243
transform 1 0 1180 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1524952243
transform 1 0 1228 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_57
timestamp 1524952243
transform 1 0 1180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1524952243
transform 1 0 1220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1524952243
transform 1 0 1228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1524952243
transform 1 0 1140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_115
timestamp 1524952243
transform 1 0 1140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1524952243
transform 1 0 1252 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1524952243
transform 1 0 1276 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1524952243
transform 1 0 1236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1524952243
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1524952243
transform 1 0 1276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1524952243
transform 1 0 1244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1524952243
transform 1 0 1252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1524952243
transform 1 0 1268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1524952243
transform 1 0 1276 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_116
timestamp 1524952243
transform 1 0 1276 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1524952243
transform 1 0 1268 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1524952243
transform 1 0 1300 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1524952243
transform 1 0 1340 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1524952243
transform 1 0 1348 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1524952243
transform 1 0 1340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1524952243
transform 1 0 1300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1524952243
transform 1 0 1324 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1524952243
transform 1 0 1372 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1524952243
transform 1 0 1364 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1524952243
transform 1 0 1348 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_63
timestamp 1524952243
transform 1 0 1356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1524952243
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1524952243
transform 1 0 1372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1524952243
transform 1 0 1332 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_117
timestamp 1524952243
transform 1 0 1348 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1524952243
transform 1 0 1420 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1524952243
transform 1 0 1388 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1524952243
transform 1 0 1428 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1524952243
transform 1 0 1428 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1524952243
transform 1 0 1396 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1524952243
transform 1 0 1404 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1524952243
transform 1 0 1412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1524952243
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1524952243
transform 1 0 1396 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1524952243
transform 1 0 1404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1524952243
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1524952243
transform 1 0 1428 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_128
timestamp 1524952243
transform 1 0 1396 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1524952243
transform 1 0 1508 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1524952243
transform 1 0 1444 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1524952243
transform 1 0 1484 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1524952243
transform 1 0 1556 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_68
timestamp 1524952243
transform 1 0 1444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1524952243
transform 1 0 1484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1524952243
transform 1 0 1540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1524952243
transform 1 0 1596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1524952243
transform 1 0 1460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1524952243
transform 1 0 1484 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1524952243
transform 1 0 1508 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1524952243
transform 1 0 1532 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1524952243
transform 1 0 1460 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1524952243
transform 1 0 1652 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1524952243
transform 1 0 1660 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_81
timestamp 1524952243
transform 1 0 1668 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1524952243
transform 1 0 1692 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1524952243
transform 1 0 1740 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_73
timestamp 1524952243
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1524952243
transform 1 0 1692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1524952243
transform 1 0 1700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1524952243
transform 1 0 1740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1524952243
transform 1 0 1556 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1524952243
transform 1 0 1596 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1524952243
transform 1 0 1644 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1524952243
transform 1 0 1764 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1524952243
transform 1 0 1820 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1524952243
transform 1 0 1836 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1524952243
transform 1 0 1796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1524952243
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1524952243
transform 1 0 1668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1524952243
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_119
timestamp 1524952243
transform 1 0 1556 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1524952243
transform 1 0 1700 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1524952243
transform 1 0 1748 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_130
timestamp 1524952243
transform 1 0 1780 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_83
timestamp 1524952243
transform 1 0 1804 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_78
timestamp 1524952243
transform 1 0 1812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1524952243
transform 1 0 1836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1524952243
transform 1 0 1804 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1524952243
transform 1 0 1820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1524952243
transform 1 0 1828 0 1 1805
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_1
timestamp 1524952243
transform 1 0 1994 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_71
timestamp 1524952243
transform 1 0 1940 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_80
timestamp 1524952243
transform 1 0 1844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1524952243
transform 1 0 1884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1524952243
transform 1 0 1940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1524952243
transform 1 0 1860 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_120
timestamp 1524952243
transform 1 0 1860 0 1 1795
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_2
timestamp 1524952243
transform 1 0 48 0 1 1770
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_0
timestamp 1524952243
transform -1 0 168 0 1 1770
box -8 -3 104 105
use NAND2X1  NAND2X1_0
timestamp 1524952243
transform 1 0 168 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_0
timestamp 1524952243
transform -1 0 208 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_0
timestamp 1524952243
transform -1 0 240 0 1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_0
timestamp 1524952243
transform -1 0 272 0 1 1770
box -8 -3 40 105
use INVX2  INVX2_1
timestamp 1524952243
transform -1 0 288 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_129
timestamp 1524952243
transform 1 0 324 0 1 1775
box -3 -3 3 3
use NAND2X1  NAND2X1_1
timestamp 1524952243
transform 1 0 288 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_2
timestamp 1524952243
transform -1 0 328 0 1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_1
timestamp 1524952243
transform 1 0 328 0 1 1770
box -8 -3 40 105
use DFFPOSX1  DFFPOSX1_1
timestamp 1524952243
transform -1 0 456 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_130
timestamp 1524952243
transform 1 0 476 0 1 1775
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_2
timestamp 1524952243
transform 1 0 456 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_131
timestamp 1524952243
transform 1 0 564 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_3
timestamp 1524952243
transform 1 0 552 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_132
timestamp 1524952243
transform 1 0 588 0 1 1775
box -3 -3 3 3
use NOR2X1  NOR2X1_0
timestamp 1524952243
transform 1 0 568 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_4
timestamp 1524952243
transform 1 0 592 0 1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_0
timestamp 1524952243
transform 1 0 608 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_5
timestamp 1524952243
transform 1 0 648 0 1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_1
timestamp 1524952243
transform -1 0 688 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_6
timestamp 1524952243
transform 1 0 688 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_1
timestamp 1524952243
transform 1 0 704 0 1 1770
box -8 -3 34 105
use INVX2  INVX2_7
timestamp 1524952243
transform 1 0 736 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_2
timestamp 1524952243
transform -1 0 784 0 1 1770
box -8 -3 34 105
use M3_M2  M3_M2_133
timestamp 1524952243
transform 1 0 796 0 1 1775
box -3 -3 3 3
use NAND3X1  NAND3X1_2
timestamp 1524952243
transform -1 0 816 0 1 1770
box -8 -3 40 105
use M3_M2  M3_M2_134
timestamp 1524952243
transform 1 0 828 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_8
timestamp 1524952243
transform -1 0 832 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_135
timestamp 1524952243
transform 1 0 868 0 1 1775
box -3 -3 3 3
use OAI21X1  OAI21X1_3
timestamp 1524952243
transform -1 0 864 0 1 1770
box -8 -3 34 105
use NOR2X1  NOR2X1_2
timestamp 1524952243
transform 1 0 864 0 1 1770
box -8 -3 32 105
use NAND3X1  NAND3X1_3
timestamp 1524952243
transform 1 0 888 0 1 1770
box -8 -3 40 105
use INVX2  INVX2_9
timestamp 1524952243
transform 1 0 920 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_4
timestamp 1524952243
transform -1 0 968 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1524952243
transform 1 0 968 0 1 1770
box -8 -3 34 105
use OR2X1  OR2X1_0
timestamp 1524952243
transform 1 0 1000 0 1 1770
box -8 -3 40 105
use DFFPOSX1  DFFPOSX1_3
timestamp 1524952243
transform -1 0 1128 0 1 1770
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_4
timestamp 1524952243
transform 1 0 1128 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_10
timestamp 1524952243
transform -1 0 1240 0 1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_1
timestamp 1524952243
transform -1 0 1280 0 1 1770
box -8 -3 46 105
use NOR2X1  NOR2X1_3
timestamp 1524952243
transform 1 0 1280 0 1 1770
box -8 -3 32 105
use OR2X1  OR2X1_1
timestamp 1524952243
transform -1 0 1336 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1524952243
transform -1 0 1368 0 1 1770
box -8 -3 40 105
use NOR2X1  NOR2X1_4
timestamp 1524952243
transform -1 0 1392 0 1 1770
box -8 -3 32 105
use AOI22X1  AOI22X1_2
timestamp 1524952243
transform 1 0 1392 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_11
timestamp 1524952243
transform 1 0 1432 0 1 1770
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_5
timestamp 1524952243
transform 1 0 1448 0 1 1770
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_6
timestamp 1524952243
transform 1 0 1544 0 1 1770
box -8 -3 104 105
use AOI22X1  AOI22X1_3
timestamp 1524952243
transform -1 0 1680 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_12
timestamp 1524952243
transform 1 0 1680 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_136
timestamp 1524952243
transform 1 0 1780 0 1 1775
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_7
timestamp 1524952243
transform -1 0 1792 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_137
timestamp 1524952243
transform 1 0 1804 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_4
timestamp 1524952243
transform 1 0 1792 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_13
timestamp 1524952243
transform 1 0 1832 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_138
timestamp 1524952243
transform 1 0 1868 0 1 1775
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_8
timestamp 1524952243
transform 1 0 1848 0 1 1770
box -8 -3 104 105
use top_module_VIA0  top_module_VIA0_3
timestamp 1524952243
transform 1 0 1970 0 1 1770
box -10 -3 10 3
use M3_M2  M3_M2_163
timestamp 1524952243
transform 1 0 132 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1524952243
transform 1 0 68 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1524952243
transform 1 0 188 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1524952243
transform 1 0 156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1524952243
transform 1 0 172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1524952243
transform 1 0 68 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1524952243
transform 1 0 132 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_185
timestamp 1524952243
transform 1 0 180 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_148
timestamp 1524952243
transform 1 0 188 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_147
timestamp 1524952243
transform 1 0 236 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1524952243
transform 1 0 212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1524952243
transform 1 0 188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1524952243
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1524952243
transform 1 0 188 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1524952243
transform 1 0 188 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1524952243
transform 1 0 252 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1524952243
transform 1 0 252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1524952243
transform 1 0 236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1524952243
transform 1 0 260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_198
timestamp 1524952243
transform 1 0 268 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1524952243
transform 1 0 308 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1524952243
transform 1 0 332 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1524952243
transform 1 0 388 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1524952243
transform 1 0 300 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_140
timestamp 1524952243
transform 1 0 300 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1524952243
transform 1 0 300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1524952243
transform 1 0 308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1524952243
transform 1 0 276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1524952243
transform 1 0 220 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1524952243
transform 1 0 236 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1524952243
transform 1 0 244 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1524952243
transform 1 0 268 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1524952243
transform 1 0 228 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1524952243
transform 1 0 236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1524952243
transform 1 0 228 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1524952243
transform 1 0 300 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_250
timestamp 1524952243
transform 1 0 292 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1524952243
transform 1 0 284 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1524952243
transform 1 0 292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1524952243
transform 1 0 404 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1524952243
transform 1 0 444 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1524952243
transform 1 0 476 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1524952243
transform 1 0 428 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_191
timestamp 1524952243
transform 1 0 340 0 1 1733
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1524952243
transform 1 0 420 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1524952243
transform 1 0 484 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1524952243
transform 1 0 516 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1524952243
transform 1 0 428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1524952243
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1524952243
transform 1 0 484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1524952243
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1524952243
transform 1 0 364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1524952243
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1524952243
transform 1 0 324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1524952243
transform 1 0 404 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1524952243
transform 1 0 356 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1524952243
transform 1 0 492 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1524952243
transform 1 0 564 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1524952243
transform 1 0 556 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1524952243
transform 1 0 580 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1524952243
transform 1 0 508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1524952243
transform 1 0 516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1524952243
transform 1 0 532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1524952243
transform 1 0 548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1524952243
transform 1 0 556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1524952243
transform 1 0 484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1524952243
transform 1 0 484 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_227
timestamp 1524952243
transform 1 0 452 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1524952243
transform 1 0 484 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1524952243
transform 1 0 420 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1524952243
transform 1 0 508 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1524952243
transform 1 0 516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1524952243
transform 1 0 524 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_201
timestamp 1524952243
transform 1 0 532 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_206
timestamp 1524952243
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1524952243
transform 1 0 556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1524952243
transform 1 0 572 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1524952243
transform 1 0 516 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1524952243
transform 1 0 524 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1524952243
transform 1 0 532 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1524952243
transform 1 0 612 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_141
timestamp 1524952243
transform 1 0 612 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1524952243
transform 1 0 620 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1524952243
transform 1 0 644 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_161
timestamp 1524952243
transform 1 0 580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1524952243
transform 1 0 604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1524952243
transform 1 0 612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1524952243
transform 1 0 620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1524952243
transform 1 0 580 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1524952243
transform 1 0 580 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1524952243
transform 1 0 572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1524952243
transform 1 0 564 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1524952243
transform 1 0 588 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1524952243
transform 1 0 628 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1524952243
transform 1 0 684 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1524952243
transform 1 0 668 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_142
timestamp 1524952243
transform 1 0 684 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1524952243
transform 1 0 700 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1524952243
transform 1 0 644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1524952243
transform 1 0 628 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1524952243
transform 1 0 612 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1524952243
transform 1 0 660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1524952243
transform 1 0 676 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1524952243
transform 1 0 700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1524952243
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1524952243
transform 1 0 668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1524952243
transform 1 0 684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1524952243
transform 1 0 644 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1524952243
transform 1 0 652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1524952243
transform 1 0 676 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1524952243
transform 1 0 644 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1524952243
transform 1 0 684 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_268
timestamp 1524952243
transform 1 0 660 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1524952243
transform 1 0 660 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_213
timestamp 1524952243
transform 1 0 708 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1524952243
transform 1 0 692 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1524952243
transform 1 0 724 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1524952243
transform 1 0 724 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1524952243
transform 1 0 764 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1524952243
transform 1 0 764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1524952243
transform 1 0 724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1524952243
transform 1 0 740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1524952243
transform 1 0 764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1524952243
transform 1 0 732 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1524952243
transform 1 0 756 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_213
timestamp 1524952243
transform 1 0 764 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1524952243
transform 1 0 740 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_269
timestamp 1524952243
transform 1 0 748 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1524952243
transform 1 0 724 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1524952243
transform 1 0 796 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1524952243
transform 1 0 812 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1524952243
transform 1 0 788 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1524952243
transform 1 0 788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1524952243
transform 1 0 796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1524952243
transform 1 0 812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1524952243
transform 1 0 788 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1524952243
transform 1 0 804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_157
timestamp 1524952243
transform 1 0 836 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1524952243
transform 1 0 860 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1524952243
transform 1 0 836 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1524952243
transform 1 0 860 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1524952243
transform 1 0 892 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1524952243
transform 1 0 860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1524952243
transform 1 0 876 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_192
timestamp 1524952243
transform 1 0 884 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1524952243
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_202
timestamp 1524952243
transform 1 0 860 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1524952243
transform 1 0 876 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1524952243
transform 1 0 884 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_214
timestamp 1524952243
transform 1 0 860 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1524952243
transform 1 0 884 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1524952243
transform 1 0 940 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1524952243
transform 1 0 940 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1524952243
transform 1 0 908 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_193
timestamp 1524952243
transform 1 0 916 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1524952243
transform 1 0 916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1524952243
transform 1 0 948 0 1 1733
box -2 -2 2 2
use M3_M2  M3_M2_177
timestamp 1524952243
transform 1 0 972 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1524952243
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1524952243
transform 1 0 980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1524952243
transform 1 0 964 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1524952243
transform 1 0 964 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1524952243
transform 1 0 1004 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1524952243
transform 1 0 996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1524952243
transform 1 0 996 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_144
timestamp 1524952243
transform 1 0 1036 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1524952243
transform 1 0 1132 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1524952243
transform 1 0 1092 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1524952243
transform 1 0 1116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1524952243
transform 1 0 1036 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1524952243
transform 1 0 1076 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1524952243
transform 1 0 1156 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1524952243
transform 1 0 1116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1524952243
transform 1 0 1132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1524952243
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1524952243
transform 1 0 1036 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1524952243
transform 1 0 1020 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1524952243
transform 1 0 1068 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_225
timestamp 1524952243
transform 1 0 1076 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_205
timestamp 1524952243
transform 1 0 1116 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_258
timestamp 1524952243
transform 1 0 1028 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1524952243
transform 1 0 1076 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_180
timestamp 1524952243
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1524952243
transform 1 0 1276 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1524952243
transform 1 0 1324 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1524952243
transform 1 0 1140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1524952243
transform 1 0 1196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1524952243
transform 1 0 1236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1524952243
transform 1 0 1244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1524952243
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_218
timestamp 1524952243
transform 1 0 1196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1524952243
transform 1 0 1244 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1524952243
transform 1 0 1140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1524952243
transform 1 0 1260 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1524952243
transform 1 0 1260 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1524952243
transform 1 0 1356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1524952243
transform 1 0 1364 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1524952243
transform 1 0 1388 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1524952243
transform 1 0 1348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1524952243
transform 1 0 1364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1524952243
transform 1 0 1524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1524952243
transform 1 0 1532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1524952243
transform 1 0 1348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1524952243
transform 1 0 1388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1524952243
transform 1 0 1444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1524952243
transform 1 0 1316 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1524952243
transform 1 0 1348 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1524952243
transform 1 0 1348 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1524952243
transform 1 0 1540 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_234
timestamp 1524952243
transform 1 0 1532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1524952243
transform 1 0 1540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1524952243
transform 1 0 1452 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_220
timestamp 1524952243
transform 1 0 1460 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1524952243
transform 1 0 1492 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_221
timestamp 1524952243
transform 1 0 1500 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1524952243
transform 1 0 1492 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1524952243
transform 1 0 1452 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1524952243
transform 1 0 1356 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1524952243
transform 1 0 1604 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1524952243
transform 1 0 1636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1524952243
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1524952243
transform 1 0 1628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1524952243
transform 1 0 1556 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1524952243
transform 1 0 1604 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1524952243
transform 1 0 1636 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1524952243
transform 1 0 1644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1524952243
transform 1 0 1660 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1524952243
transform 1 0 1628 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1524952243
transform 1 0 1660 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1524952243
transform 1 0 1756 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1524952243
transform 1 0 1716 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_186
timestamp 1524952243
transform 1 0 1748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1524952243
transform 1 0 1756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1524952243
transform 1 0 1780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1524952243
transform 1 0 1868 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1524952243
transform 1 0 1748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1524952243
transform 1 0 1716 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1524952243
transform 1 0 1740 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1524952243
transform 1 0 1788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1524952243
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1524952243
transform 1 0 1884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1524952243
transform 1 0 1900 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1524952243
transform 1 0 1788 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1524952243
transform 1 0 1868 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1524952243
transform 1 0 1772 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1524952243
transform 1 0 1900 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1524952243
transform 1 0 1932 0 1 1735
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_4
timestamp 1524952243
transform 1 0 24 0 1 1670
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_9
timestamp 1524952243
transform -1 0 168 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_14
timestamp 1524952243
transform 1 0 168 0 -1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_6
timestamp 1524952243
transform -1 0 216 0 -1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_5
timestamp 1524952243
transform -1 0 248 0 -1 1770
box -8 -3 40 105
use INVX2  INVX2_15
timestamp 1524952243
transform 1 0 248 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_6
timestamp 1524952243
transform 1 0 264 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1524952243
transform 1 0 296 0 -1 1770
box -8 -3 40 105
use DFFPOSX1  DFFPOSX1_10
timestamp 1524952243
transform 1 0 328 0 -1 1770
box -8 -3 104 105
use XOR2X1  XOR2X1_0
timestamp 1524952243
transform 1 0 424 0 -1 1770
box -8 -3 64 105
use OAI21X1  OAI21X1_7
timestamp 1524952243
transform -1 0 512 0 -1 1770
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1524952243
transform 1 0 512 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_16
timestamp 1524952243
transform 1 0 552 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1524952243
transform -1 0 584 0 -1 1770
box -9 -3 26 105
use OR2X1  OR2X1_3
timestamp 1524952243
transform -1 0 616 0 -1 1770
box -8 -3 40 105
use OAI21X1  OAI21X1_8
timestamp 1524952243
transform 1 0 616 0 -1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_7
timestamp 1524952243
transform -1 0 680 0 -1 1770
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1524952243
transform -1 0 712 0 -1 1770
box -7 -3 39 105
use INVX2  INVX2_18
timestamp 1524952243
transform 1 0 712 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_8
timestamp 1524952243
transform 1 0 728 0 -1 1770
box -8 -3 40 105
use OAI21X1  OAI21X1_9
timestamp 1524952243
transform 1 0 760 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_19
timestamp 1524952243
transform 1 0 792 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1524952243
transform 1 0 808 0 -1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_10
timestamp 1524952243
transform 1 0 824 0 -1 1770
box -8 -3 34 105
use AOI21X1  AOI21X1_1
timestamp 1524952243
transform -1 0 888 0 -1 1770
box -7 -3 39 105
use NOR2X1  NOR2X1_5
timestamp 1524952243
transform 1 0 888 0 -1 1770
box -8 -3 32 105
use AOI21X1  AOI21X1_2
timestamp 1524952243
transform 1 0 912 0 -1 1770
box -7 -3 39 105
use OAI21X1  OAI21X1_11
timestamp 1524952243
transform -1 0 976 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_21
timestamp 1524952243
transform 1 0 976 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1524952243
transform 1 0 992 0 -1 1770
box -9 -3 26 105
use NAND2X1  NAND2X1_2
timestamp 1524952243
transform 1 0 1008 0 -1 1770
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_11
timestamp 1524952243
transform -1 0 1128 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_23
timestamp 1524952243
transform 1 0 1128 0 -1 1770
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_12
timestamp 1524952243
transform 1 0 1144 0 -1 1770
box -8 -3 104 105
use AND2X2  AND2X2_0
timestamp 1524952243
transform -1 0 1272 0 -1 1770
box -8 -3 40 105
use HAX1  HAX1_0
timestamp 1524952243
transform -1 0 1352 0 -1 1770
box -5 -3 84 105
use DFFPOSX1  DFFPOSX1_13
timestamp 1524952243
transform 1 0 1352 0 -1 1770
box -8 -3 104 105
use HAX1  HAX1_1
timestamp 1524952243
transform -1 0 1528 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1524952243
transform 1 0 1528 0 -1 1770
box -5 -3 84 105
use AND2X2  AND2X2_1
timestamp 1524952243
transform -1 0 1640 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1524952243
transform -1 0 1672 0 -1 1770
box -8 -3 40 105
use M3_M2  M3_M2_256
timestamp 1524952243
transform 1 0 1748 0 1 1675
box -3 -3 3 3
use HAX1  HAX1_3
timestamp 1524952243
transform -1 0 1752 0 -1 1770
box -5 -3 84 105
use OAI21X1  OAI21X1_12
timestamp 1524952243
transform -1 0 1784 0 -1 1770
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_14
timestamp 1524952243
transform -1 0 1880 0 -1 1770
box -8 -3 104 105
use M3_M2  M3_M2_257
timestamp 1524952243
transform 1 0 1892 0 1 1675
box -3 -3 3 3
use AND2X2  AND2X2_3
timestamp 1524952243
transform -1 0 1912 0 -1 1770
box -8 -3 40 105
use FILL  FILL_0
timestamp 1524952243
transform 1 0 1912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1
timestamp 1524952243
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2
timestamp 1524952243
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3
timestamp 1524952243
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_5
timestamp 1524952243
transform 1 0 1994 0 1 1670
box -10 -3 10 3
use M3_M2  M3_M2_276
timestamp 1524952243
transform 1 0 132 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1524952243
transform 1 0 172 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1524952243
transform 1 0 252 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1524952243
transform 1 0 284 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1524952243
transform 1 0 268 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_270
timestamp 1524952243
transform 1 0 300 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1524952243
transform 1 0 284 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1524952243
transform 1 0 68 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1524952243
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1524952243
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1524952243
transform 1 0 156 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1524952243
transform 1 0 180 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_285
timestamp 1524952243
transform 1 0 188 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1524952243
transform 1 0 228 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_286
timestamp 1524952243
transform 1 0 244 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_300
timestamp 1524952243
transform 1 0 252 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_347
timestamp 1524952243
transform 1 0 180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1524952243
transform 1 0 268 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_321
timestamp 1524952243
transform 1 0 156 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1524952243
transform 1 0 268 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1524952243
transform 1 0 308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1524952243
transform 1 0 292 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1524952243
transform 1 0 308 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1524952243
transform 1 0 340 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_288
timestamp 1524952243
transform 1 0 316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1524952243
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_311
timestamp 1524952243
transform 1 0 324 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_349
timestamp 1524952243
transform 1 0 332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1524952243
transform 1 0 348 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_302
timestamp 1524952243
transform 1 0 348 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_290
timestamp 1524952243
transform 1 0 356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1524952243
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1524952243
transform 1 0 404 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1524952243
transform 1 0 404 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1524952243
transform 1 0 428 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1524952243
transform 1 0 420 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1524952243
transform 1 0 412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1524952243
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_278
timestamp 1524952243
transform 1 0 468 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1524952243
transform 1 0 508 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_293
timestamp 1524952243
transform 1 0 460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1524952243
transform 1 0 468 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_304
timestamp 1524952243
transform 1 0 484 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1524952243
transform 1 0 628 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1524952243
transform 1 0 676 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_276
timestamp 1524952243
transform 1 0 684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1524952243
transform 1 0 508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1524952243
transform 1 0 564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1524952243
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1524952243
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1524952243
transform 1 0 668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1524952243
transform 1 0 676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1524952243
transform 1 0 452 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1524952243
transform 1 0 444 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_343
timestamp 1524952243
transform 1 0 484 0 1 1607
box -2 -2 2 2
use M3_M2  M3_M2_335
timestamp 1524952243
transform 1 0 484 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_352
timestamp 1524952243
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1524952243
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1524952243
transform 1 0 732 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1524952243
transform 1 0 740 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1524952243
transform 1 0 804 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1524952243
transform 1 0 700 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1524952243
transform 1 0 804 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1524952243
transform 1 0 716 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_301
timestamp 1524952243
transform 1 0 740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1524952243
transform 1 0 796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1524952243
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1524952243
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1524952243
transform 1 0 716 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1524952243
transform 1 0 740 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1524952243
transform 1 0 836 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_304
timestamp 1524952243
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1524952243
transform 1 0 820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1524952243
transform 1 0 804 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_336
timestamp 1524952243
transform 1 0 716 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1524952243
transform 1 0 732 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1524952243
transform 1 0 804 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1524952243
transform 1 0 852 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_305
timestamp 1524952243
transform 1 0 844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1524952243
transform 1 0 852 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_285
timestamp 1524952243
transform 1 0 868 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_307
timestamp 1524952243
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1524952243
transform 1 0 860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1524952243
transform 1 0 868 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1524952243
transform 1 0 900 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_308
timestamp 1524952243
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1524952243
transform 1 0 908 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_313
timestamp 1524952243
transform 1 0 900 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1524952243
transform 1 0 900 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1524952243
transform 1 0 900 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_310
timestamp 1524952243
transform 1 0 916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1524952243
transform 1 0 924 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_306
timestamp 1524952243
transform 1 0 948 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_312
timestamp 1524952243
transform 1 0 956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1524952243
transform 1 0 932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1524952243
transform 1 0 940 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1524952243
transform 1 0 932 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_313
timestamp 1524952243
transform 1 0 980 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_307
timestamp 1524952243
transform 1 0 988 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_314
timestamp 1524952243
transform 1 0 996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1524952243
transform 1 0 964 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1524952243
transform 1 0 964 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_361
timestamp 1524952243
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1524952243
transform 1 0 1004 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1524952243
transform 1 0 1036 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1524952243
transform 1 0 1028 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1524952243
transform 1 0 1020 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1524952243
transform 1 0 1068 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1524952243
transform 1 0 1052 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1524952243
transform 1 0 1108 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1524952243
transform 1 0 1156 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_315
timestamp 1524952243
transform 1 0 1036 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_308
timestamp 1524952243
transform 1 0 1044 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_362
timestamp 1524952243
transform 1 0 1028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1524952243
transform 1 0 1044 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1524952243
transform 1 0 1012 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1524952243
transform 1 0 1180 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1524952243
transform 1 0 1268 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1524952243
transform 1 0 1284 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1524952243
transform 1 0 1316 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1524952243
transform 1 0 1220 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1524952243
transform 1 0 1252 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1524952243
transform 1 0 1316 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1524952243
transform 1 0 1340 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_316
timestamp 1524952243
transform 1 0 1052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1524952243
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1524952243
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1524952243
transform 1 0 1156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1524952243
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1524952243
transform 1 0 1188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1524952243
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1524952243
transform 1 0 1068 0 1 1607
box -2 -2 2 2
use M3_M2  M3_M2_315
timestamp 1524952243
transform 1 0 1092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1524952243
transform 1 0 1052 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1524952243
transform 1 0 1100 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1524952243
transform 1 0 1036 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1524952243
transform 1 0 1164 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_364
timestamp 1524952243
transform 1 0 1172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1524952243
transform 1 0 1180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1524952243
transform 1 0 1196 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_309
timestamp 1524952243
transform 1 0 1252 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1524952243
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1524952243
transform 1 0 1292 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1524952243
transform 1 0 1316 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_317
timestamp 1524952243
transform 1 0 1276 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1524952243
transform 1 0 1388 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1524952243
transform 1 0 1380 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1524952243
transform 1 0 1420 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_325
timestamp 1524952243
transform 1 0 1356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1524952243
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1524952243
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1524952243
transform 1 0 1396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1524952243
transform 1 0 1412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1524952243
transform 1 0 1420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1524952243
transform 1 0 1476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1524952243
transform 1 0 1284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1524952243
transform 1 0 1292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1524952243
transform 1 0 1340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1524952243
transform 1 0 1348 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_326
timestamp 1524952243
transform 1 0 1340 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1524952243
transform 1 0 1388 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_318
timestamp 1524952243
transform 1 0 1396 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_372
timestamp 1524952243
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_319
timestamp 1524952243
transform 1 0 1468 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_345
timestamp 1524952243
transform 1 0 1500 0 1 1607
box -2 -2 2 2
use M3_M2  M3_M2_327
timestamp 1524952243
transform 1 0 1500 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1524952243
transform 1 0 1412 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1524952243
transform 1 0 1460 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1524952243
transform 1 0 1564 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1524952243
transform 1 0 1612 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1524952243
transform 1 0 1708 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1524952243
transform 1 0 1756 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_332
timestamp 1524952243
transform 1 0 1564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1524952243
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1524952243
transform 1 0 1620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1524952243
transform 1 0 1636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1524952243
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1524952243
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1524952243
transform 1 0 1748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1524952243
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1524952243
transform 1 0 1772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1524952243
transform 1 0 1524 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1524952243
transform 1 0 1564 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1524952243
transform 1 0 1524 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1524952243
transform 1 0 1572 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_374
timestamp 1524952243
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1524952243
transform 1 0 1628 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1524952243
transform 1 0 1620 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_376
timestamp 1524952243
transform 1 0 1668 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_348
timestamp 1524952243
transform 1 0 1668 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_279
timestamp 1524952243
transform 1 0 1836 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1524952243
transform 1 0 1892 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1524952243
transform 1 0 1932 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1524952243
transform 1 0 1852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1524952243
transform 1 0 1860 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1524952243
transform 1 0 1852 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1524952243
transform 1 0 1860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1524952243
transform 1 0 1868 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1524952243
transform 1 0 1764 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1524952243
transform 1 0 1780 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1524952243
transform 1 0 1828 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1524952243
transform 1 0 1860 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1524952243
transform 1 0 1940 0 1 1595
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_6
timestamp 1524952243
transform 1 0 48 0 1 1570
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_15
timestamp 1524952243
transform -1 0 168 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_24
timestamp 1524952243
transform -1 0 184 0 1 1570
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_16
timestamp 1524952243
transform -1 0 280 0 1 1570
box -8 -3 104 105
use NAND3X1  NAND3X1_9
timestamp 1524952243
transform 1 0 280 0 1 1570
box -8 -3 40 105
use INVX2  INVX2_25
timestamp 1524952243
transform -1 0 328 0 1 1570
box -9 -3 26 105
use NAND2X1  NAND2X1_3
timestamp 1524952243
transform 1 0 328 0 1 1570
box -8 -3 32 105
use INVX2  INVX2_26
timestamp 1524952243
transform 1 0 352 0 1 1570
box -9 -3 26 105
use FILL  FILL_4
timestamp 1524952243
transform 1 0 368 0 1 1570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1524952243
transform 1 0 376 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1524952243
transform -1 0 408 0 1 1570
box -8 -3 32 105
use FILL  FILL_6
timestamp 1524952243
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1524952243
transform 1 0 416 0 1 1570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1524952243
transform 1 0 424 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_349
timestamp 1524952243
transform 1 0 460 0 1 1575
box -3 -3 3 3
use NAND2X1  NAND2X1_5
timestamp 1524952243
transform -1 0 456 0 1 1570
box -8 -3 32 105
use INVX2  INVX2_27
timestamp 1524952243
transform 1 0 456 0 1 1570
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_17
timestamp 1524952243
transform 1 0 472 0 1 1570
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_18
timestamp 1524952243
transform -1 0 664 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_28
timestamp 1524952243
transform -1 0 680 0 1 1570
box -9 -3 26 105
use NAND2X1  NAND2X1_6
timestamp 1524952243
transform -1 0 704 0 1 1570
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_19
timestamp 1524952243
transform 1 0 704 0 1 1570
box -8 -3 104 105
use AOI21X1  AOI21X1_3
timestamp 1524952243
transform -1 0 832 0 1 1570
box -7 -3 39 105
use INVX2  INVX2_29
timestamp 1524952243
transform 1 0 832 0 1 1570
box -9 -3 26 105
use NOR2X1  NOR2X1_6
timestamp 1524952243
transform -1 0 872 0 1 1570
box -8 -3 32 105
use AOI21X1  AOI21X1_4
timestamp 1524952243
transform 1 0 872 0 1 1570
box -7 -3 39 105
use INVX2  INVX2_30
timestamp 1524952243
transform -1 0 920 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1524952243
transform -1 0 936 0 1 1570
box -9 -3 26 105
use BUFX2  BUFX2_0
timestamp 1524952243
transform -1 0 960 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1524952243
transform -1 0 984 0 1 1570
box -5 -3 28 105
use INVX2  INVX2_32
timestamp 1524952243
transform -1 0 1000 0 1 1570
box -9 -3 26 105
use BUFX2  BUFX2_2
timestamp 1524952243
transform 1 0 1000 0 1 1570
box -5 -3 28 105
use INVX2  INVX2_33
timestamp 1524952243
transform 1 0 1024 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1524952243
transform 1 0 1040 0 1 1570
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_20
timestamp 1524952243
transform 1 0 1056 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1524952243
transform -1 0 1168 0 1 1570
box -9 -3 26 105
use M3_M2  M3_M2_350
timestamp 1524952243
transform 1 0 1196 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_5
timestamp 1524952243
transform 1 0 1168 0 1 1570
box -8 -3 46 105
use HAX1  HAX1_4
timestamp 1524952243
transform -1 0 1288 0 1 1570
box -5 -3 84 105
use XOR2X1  XOR2X1_1
timestamp 1524952243
transform 1 0 1288 0 1 1570
box -8 -3 64 105
use AND2X2  AND2X2_4
timestamp 1524952243
transform 1 0 1344 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_351
timestamp 1524952243
transform 1 0 1404 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_6
timestamp 1524952243
transform 1 0 1376 0 1 1570
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_21
timestamp 1524952243
transform -1 0 1512 0 1 1570
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_22
timestamp 1524952243
transform 1 0 1512 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_352
timestamp 1524952243
transform 1 0 1620 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_36
timestamp 1524952243
transform -1 0 1624 0 1 1570
box -9 -3 26 105
use M3_M2  M3_M2_353
timestamp 1524952243
transform 1 0 1644 0 1 1575
box -3 -3 3 3
use AND2X2  AND2X2_5
timestamp 1524952243
transform 1 0 1624 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_354
timestamp 1524952243
transform 1 0 1732 0 1 1575
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_23
timestamp 1524952243
transform 1 0 1656 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_355
timestamp 1524952243
transform 1 0 1772 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1524952243
transform 1 0 1796 0 1 1575
box -3 -3 3 3
use AND2X2  AND2X2_6
timestamp 1524952243
transform -1 0 1784 0 1 1570
box -8 -3 40 105
use HAX1  HAX1_5
timestamp 1524952243
transform -1 0 1864 0 1 1570
box -5 -3 84 105
use HAX1  HAX1_6
timestamp 1524952243
transform 1 0 1864 0 1 1570
box -5 -3 84 105
use top_module_VIA0  top_module_VIA0_7
timestamp 1524952243
transform 1 0 1970 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_387
timestamp 1524952243
transform 1 0 68 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_385
timestamp 1524952243
transform 1 0 156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1524952243
transform 1 0 68 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_398
timestamp 1524952243
transform 1 0 84 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1524952243
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_399
timestamp 1524952243
transform 1 0 156 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1524952243
transform 1 0 260 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_386
timestamp 1524952243
transform 1 0 180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1524952243
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_408
timestamp 1524952243
transform 1 0 220 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1524952243
transform 1 0 204 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1524952243
transform 1 0 284 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_382
timestamp 1524952243
transform 1 0 292 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1524952243
transform 1 0 292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1524952243
transform 1 0 276 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_400
timestamp 1524952243
transform 1 0 284 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1524952243
transform 1 0 284 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1524952243
transform 1 0 292 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1524952243
transform 1 0 284 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1524952243
transform 1 0 308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1524952243
transform 1 0 340 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1524952243
transform 1 0 324 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_388
timestamp 1524952243
transform 1 0 340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1524952243
transform 1 0 348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1524952243
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1524952243
transform 1 0 316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1524952243
transform 1 0 324 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_401
timestamp 1524952243
transform 1 0 332 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1524952243
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_402
timestamp 1524952243
transform 1 0 348 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1524952243
transform 1 0 388 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1524952243
transform 1 0 380 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_432
timestamp 1524952243
transform 1 0 372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1524952243
transform 1 0 380 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_432
timestamp 1524952243
transform 1 0 316 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_484
timestamp 1524952243
transform 1 0 340 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_410
timestamp 1524952243
transform 1 0 356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1524952243
transform 1 0 388 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1524952243
transform 1 0 444 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1524952243
transform 1 0 484 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1524952243
transform 1 0 428 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1524952243
transform 1 0 468 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_390
timestamp 1524952243
transform 1 0 428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1524952243
transform 1 0 444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1524952243
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1524952243
transform 1 0 396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1524952243
transform 1 0 404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1524952243
transform 1 0 412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1524952243
transform 1 0 364 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_433
timestamp 1524952243
transform 1 0 372 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1524952243
transform 1 0 340 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1524952243
transform 1 0 356 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1524952243
transform 1 0 396 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_411
timestamp 1524952243
transform 1 0 404 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_437
timestamp 1524952243
transform 1 0 468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1524952243
transform 1 0 524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1524952243
transform 1 0 532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1524952243
transform 1 0 428 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_434
timestamp 1524952243
transform 1 0 396 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1524952243
transform 1 0 476 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_393
timestamp 1524952243
transform 1 0 556 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_357
timestamp 1524952243
transform 1 0 660 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1524952243
transform 1 0 580 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1524952243
transform 1 0 668 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1524952243
transform 1 0 684 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_394
timestamp 1524952243
transform 1 0 580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1524952243
transform 1 0 596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1524952243
transform 1 0 684 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1524952243
transform 1 0 572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1524952243
transform 1 0 548 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_435
timestamp 1524952243
transform 1 0 532 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1524952243
transform 1 0 524 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1524952243
transform 1 0 556 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1524952243
transform 1 0 564 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_441
timestamp 1524952243
transform 1 0 620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1524952243
transform 1 0 676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1524952243
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1524952243
transform 1 0 620 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1524952243
transform 1 0 628 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1524952243
transform 1 0 684 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1524952243
transform 1 0 644 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_383
timestamp 1524952243
transform 1 0 716 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1524952243
transform 1 0 716 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1524952243
transform 1 0 820 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1524952243
transform 1 0 908 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1524952243
transform 1 0 732 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1524952243
transform 1 0 748 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1524952243
transform 1 0 836 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_397
timestamp 1524952243
transform 1 0 732 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_391
timestamp 1524952243
transform 1 0 740 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_398
timestamp 1524952243
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_367
timestamp 1524952243
transform 1 0 956 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_399
timestamp 1524952243
transform 1 0 916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1524952243
transform 1 0 932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1524952243
transform 1 0 740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1524952243
transform 1 0 780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1524952243
transform 1 0 836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1524952243
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1524952243
transform 1 0 932 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1524952243
transform 1 0 732 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1524952243
transform 1 0 780 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1524952243
transform 1 0 724 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1524952243
transform 1 0 828 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_401
timestamp 1524952243
transform 1 0 956 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_392
timestamp 1524952243
transform 1 0 996 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_402
timestamp 1524952243
transform 1 0 1044 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_393
timestamp 1524952243
transform 1 0 1052 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_403
timestamp 1524952243
transform 1 0 1060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1524952243
transform 1 0 1084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1524952243
transform 1 0 1092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1524952243
transform 1 0 980 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_404
timestamp 1524952243
transform 1 0 1020 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_450
timestamp 1524952243
transform 1 0 1036 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1524952243
transform 1 0 1044 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1524952243
transform 1 0 932 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1524952243
transform 1 0 956 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1524952243
transform 1 0 980 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1524952243
transform 1 0 1028 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1524952243
transform 1 0 1100 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1524952243
transform 1 0 1292 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1524952243
transform 1 0 1220 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_406
timestamp 1524952243
transform 1 0 1124 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_395
timestamp 1524952243
transform 1 0 1204 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_407
timestamp 1524952243
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_384
timestamp 1524952243
transform 1 0 1332 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_408
timestamp 1524952243
transform 1 0 1332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1524952243
transform 1 0 1340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1524952243
transform 1 0 1052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1524952243
transform 1 0 1060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1524952243
transform 1 0 1076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1524952243
transform 1 0 1100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1524952243
transform 1 0 1108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1524952243
transform 1 0 1148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1524952243
transform 1 0 1204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1524952243
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1524952243
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1524952243
transform 1 0 1308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1524952243
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_419
timestamp 1524952243
transform 1 0 1108 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1524952243
transform 1 0 1148 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1524952243
transform 1 0 1124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1524952243
transform 1 0 1268 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1524952243
transform 1 0 1308 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1524952243
transform 1 0 1380 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1524952243
transform 1 0 1380 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_410
timestamp 1524952243
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1524952243
transform 1 0 1468 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_359
timestamp 1524952243
transform 1 0 1564 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_412
timestamp 1524952243
transform 1 0 1564 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_370
timestamp 1524952243
transform 1 0 1604 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1524952243
transform 1 0 1628 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_413
timestamp 1524952243
transform 1 0 1596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1524952243
transform 1 0 1604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1524952243
transform 1 0 1620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1524952243
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1524952243
transform 1 0 1364 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1524952243
transform 1 0 1404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1524952243
transform 1 0 1460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1524952243
transform 1 0 1476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1524952243
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1524952243
transform 1 0 1540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1524952243
transform 1 0 1580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1524952243
transform 1 0 1588 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_423
timestamp 1524952243
transform 1 0 1364 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1524952243
transform 1 0 1404 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1524952243
transform 1 0 1540 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1524952243
transform 1 0 1580 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1524952243
transform 1 0 1484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1524952243
transform 1 0 1604 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1524952243
transform 1 0 1644 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_416
timestamp 1524952243
transform 1 0 1644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1524952243
transform 1 0 1732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1524952243
transform 1 0 1612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1524952243
transform 1 0 1628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1524952243
transform 1 0 1668 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_444
timestamp 1524952243
transform 1 0 1588 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1524952243
transform 1 0 1748 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1524952243
transform 1 0 1780 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1524952243
transform 1 0 1804 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_418
timestamp 1524952243
transform 1 0 1756 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1524952243
transform 1 0 1772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1524952243
transform 1 0 1748 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_407
timestamp 1524952243
transform 1 0 1756 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_475
timestamp 1524952243
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1524952243
transform 1 0 1772 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1524952243
transform 1 0 1756 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1524952243
transform 1 0 1772 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1524952243
transform 1 0 1788 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_420
timestamp 1524952243
transform 1 0 1796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1524952243
transform 1 0 1812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1524952243
transform 1 0 1820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1524952243
transform 1 0 1788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1524952243
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1524952243
transform 1 0 1828 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_429
timestamp 1524952243
transform 1 0 1812 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_480
timestamp 1524952243
transform 1 0 1844 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_430
timestamp 1524952243
transform 1 0 1844 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1524952243
transform 1 0 1860 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_423
timestamp 1524952243
transform 1 0 1860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1524952243
transform 1 0 1884 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1524952243
transform 1 0 1940 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_431
timestamp 1524952243
transform 1 0 1884 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1524952243
transform 1 0 1852 0 1 1505
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_8
timestamp 1524952243
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_24
timestamp 1524952243
transform -1 0 168 0 -1 1570
box -8 -3 104 105
use M3_M2  M3_M2_453
timestamp 1524952243
transform 1 0 196 0 1 1475
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_25
timestamp 1524952243
transform 1 0 168 0 -1 1570
box -8 -3 104 105
use M3_M2  M3_M2_454
timestamp 1524952243
transform 1 0 284 0 1 1475
box -3 -3 3 3
use NAND2X1  NAND2X1_7
timestamp 1524952243
transform 1 0 264 0 -1 1570
box -8 -3 32 105
use M3_M2  M3_M2_455
timestamp 1524952243
transform 1 0 316 0 1 1475
box -3 -3 3 3
use NOR2X1  NOR2X1_7
timestamp 1524952243
transform 1 0 288 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_13
timestamp 1524952243
transform 1 0 312 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_8
timestamp 1524952243
transform 1 0 344 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_14
timestamp 1524952243
transform 1 0 368 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1524952243
transform 1 0 400 0 -1 1570
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_26
timestamp 1524952243
transform 1 0 432 0 -1 1570
box -8 -3 104 105
use NAND2X1  NAND2X1_9
timestamp 1524952243
transform 1 0 528 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_16
timestamp 1524952243
transform -1 0 584 0 -1 1570
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_27
timestamp 1524952243
transform 1 0 584 0 -1 1570
box -8 -3 104 105
use AOI21X1  AOI21X1_5
timestamp 1524952243
transform 1 0 680 0 -1 1570
box -7 -3 39 105
use NOR2X1  NOR2X1_8
timestamp 1524952243
transform -1 0 736 0 -1 1570
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_28
timestamp 1524952243
transform -1 0 832 0 -1 1570
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_29
timestamp 1524952243
transform -1 0 928 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_37
timestamp 1524952243
transform 1 0 928 0 -1 1570
box -9 -3 26 105
use M3_M2  M3_M2_456
timestamp 1524952243
transform 1 0 1012 0 1 1475
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_30
timestamp 1524952243
transform 1 0 944 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_38
timestamp 1524952243
transform 1 0 1040 0 -1 1570
box -9 -3 26 105
use M3_M2  M3_M2_457
timestamp 1524952243
transform 1 0 1084 0 1 1475
box -3 -3 3 3
use AOI22X1  AOI22X1_7
timestamp 1524952243
transform -1 0 1096 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_39
timestamp 1524952243
transform 1 0 1096 0 -1 1570
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_31
timestamp 1524952243
transform 1 0 1112 0 -1 1570
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_32
timestamp 1524952243
transform -1 0 1304 0 -1 1570
box -8 -3 104 105
use AND2X2  AND2X2_7
timestamp 1524952243
transform -1 0 1336 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1524952243
transform 1 0 1336 0 -1 1570
box -8 -3 40 105
use DFFPOSX1  DFFPOSX1_33
timestamp 1524952243
transform 1 0 1368 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_40
timestamp 1524952243
transform 1 0 1464 0 -1 1570
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_34
timestamp 1524952243
transform -1 0 1576 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_41
timestamp 1524952243
transform -1 0 1592 0 -1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_8
timestamp 1524952243
transform 1 0 1592 0 -1 1570
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_35
timestamp 1524952243
transform 1 0 1632 0 -1 1570
box -8 -3 104 105
use AOI22X1  AOI22X1_9
timestamp 1524952243
transform -1 0 1768 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_42
timestamp 1524952243
transform 1 0 1768 0 -1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_10
timestamp 1524952243
transform -1 0 1824 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_43
timestamp 1524952243
transform 1 0 1824 0 -1 1570
box -9 -3 26 105
use FILL  FILL_9
timestamp 1524952243
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_36
timestamp 1524952243
transform 1 0 1848 0 -1 1570
box -8 -3 104 105
use top_module_VIA0  top_module_VIA0_9
timestamp 1524952243
transform 1 0 1994 0 1 1470
box -10 -3 10 3
use M2_M1  M2_M1_496
timestamp 1524952243
transform 1 0 76 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1524952243
transform 1 0 132 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_497
timestamp 1524952243
transform 1 0 140 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_458
timestamp 1524952243
transform 1 0 220 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_489
timestamp 1524952243
transform 1 0 220 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1524952243
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1524952243
transform 1 0 204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1524952243
transform 1 0 164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1524952243
transform 1 0 180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1524952243
transform 1 0 196 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_498
timestamp 1524952243
transform 1 0 220 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1524952243
transform 1 0 276 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1524952243
transform 1 0 308 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_490
timestamp 1524952243
transform 1 0 308 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1524952243
transform 1 0 260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1524952243
transform 1 0 284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1524952243
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1524952243
transform 1 0 340 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1524952243
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_499
timestamp 1524952243
transform 1 0 324 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1524952243
transform 1 0 380 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1524952243
transform 1 0 372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1524952243
transform 1 0 388 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1524952243
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1524952243
transform 1 0 364 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_505
timestamp 1524952243
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1524952243
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1524952243
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1524952243
transform 1 0 228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1524952243
transform 1 0 276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1524952243
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1524952243
transform 1 0 332 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1524952243
transform 1 0 348 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1524952243
transform 1 0 340 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_507
timestamp 1524952243
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1524952243
transform 1 0 380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1524952243
transform 1 0 388 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_569
timestamp 1524952243
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1524952243
transform 1 0 420 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_507
timestamp 1524952243
transform 1 0 412 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1524952243
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1524952243
transform 1 0 444 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1524952243
transform 1 0 460 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1524952243
transform 1 0 476 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_509
timestamp 1524952243
transform 1 0 428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1524952243
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_501
timestamp 1524952243
transform 1 0 452 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_511
timestamp 1524952243
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1524952243
transform 1 0 436 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_508
timestamp 1524952243
transform 1 0 444 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1524952243
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1524952243
transform 1 0 460 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1524952243
transform 1 0 524 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1524952243
transform 1 0 540 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_491
timestamp 1524952243
transform 1 0 524 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1524952243
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1524952243
transform 1 0 492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1524952243
transform 1 0 508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1524952243
transform 1 0 524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1524952243
transform 1 0 468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1524952243
transform 1 0 476 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1524952243
transform 1 0 484 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_575
timestamp 1524952243
transform 1 0 500 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1524952243
transform 1 0 428 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1524952243
transform 1 0 468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1524952243
transform 1 0 428 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1524952243
transform 1 0 500 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1524952243
transform 1 0 548 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_576
timestamp 1524952243
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1524952243
transform 1 0 548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1524952243
transform 1 0 556 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_519
timestamp 1524952243
transform 1 0 548 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1524952243
transform 1 0 572 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1524952243
transform 1 0 660 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_493
timestamp 1524952243
transform 1 0 572 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1524952243
transform 1 0 572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1524952243
transform 1 0 580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1524952243
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1524952243
transform 1 0 660 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_535
timestamp 1524952243
transform 1 0 620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1524952243
transform 1 0 644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1524952243
transform 1 0 700 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_518
timestamp 1524952243
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1524952243
transform 1 0 764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1524952243
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1524952243
transform 1 0 772 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_537
timestamp 1524952243
transform 1 0 716 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1524952243
transform 1 0 772 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1524952243
transform 1 0 820 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1524952243
transform 1 0 820 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1524952243
transform 1 0 788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1524952243
transform 1 0 804 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1524952243
transform 1 0 796 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1524952243
transform 1 0 788 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_522
timestamp 1524952243
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1524952243
transform 1 0 828 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_512
timestamp 1524952243
transform 1 0 844 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1524952243
transform 1 0 868 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1524952243
transform 1 0 932 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_523
timestamp 1524952243
transform 1 0 892 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1524952243
transform 1 0 948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1524952243
transform 1 0 956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1524952243
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1524952243
transform 1 0 868 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1524952243
transform 1 0 916 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1524952243
transform 1 0 852 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1524952243
transform 1 0 892 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1524952243
transform 1 0 948 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1524952243
transform 1 0 868 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1524952243
transform 1 0 980 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1524952243
transform 1 0 980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1524952243
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1524952243
transform 1 0 1004 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1524952243
transform 1 0 1036 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1524952243
transform 1 0 1060 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1524952243
transform 1 0 1012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1524952243
transform 1 0 1052 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1524952243
transform 1 0 1100 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1524952243
transform 1 0 1196 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_495
timestamp 1524952243
transform 1 0 1156 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1524952243
transform 1 0 1108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1524952243
transform 1 0 1116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1524952243
transform 1 0 1124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1524952243
transform 1 0 1140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1524952243
transform 1 0 972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1524952243
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1524952243
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1524952243
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1524952243
transform 1 0 1028 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_524
timestamp 1524952243
transform 1 0 988 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1524952243
transform 1 0 1052 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_589
timestamp 1524952243
transform 1 0 1132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1524952243
transform 1 0 1196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1524952243
transform 1 0 1236 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1524952243
transform 1 0 1276 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1524952243
transform 1 0 1300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1524952243
transform 1 0 1348 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1524952243
transform 1 0 1380 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1524952243
transform 1 0 1364 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1524952243
transform 1 0 1404 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1524952243
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1524952243
transform 1 0 1300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1524952243
transform 1 0 1324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1524952243
transform 1 0 1348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1524952243
transform 1 0 1364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1524952243
transform 1 0 1380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1524952243
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1524952243
transform 1 0 1404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1524952243
transform 1 0 1244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1524952243
transform 1 0 1252 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1524952243
transform 1 0 1244 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_592
timestamp 1524952243
transform 1 0 1300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1524952243
transform 1 0 1308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1524952243
transform 1 0 1332 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1524952243
transform 1 0 1348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1524952243
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1524952243
transform 1 0 1372 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1524952243
transform 1 0 1300 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1524952243
transform 1 0 1332 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1524952243
transform 1 0 1388 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1524952243
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1524952243
transform 1 0 1412 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1524952243
transform 1 0 1420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_528
timestamp 1524952243
transform 1 0 1372 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1524952243
transform 1 0 1412 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1524952243
transform 1 0 1380 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1524952243
transform 1 0 1396 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1524952243
transform 1 0 1468 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_545
timestamp 1524952243
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_466
timestamp 1524952243
transform 1 0 1564 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1524952243
transform 1 0 1532 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1524952243
transform 1 0 1604 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1524952243
transform 1 0 1636 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_546
timestamp 1524952243
transform 1 0 1532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1524952243
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1524952243
transform 1 0 1580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1524952243
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1524952243
transform 1 0 1508 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1524952243
transform 1 0 1588 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1524952243
transform 1 0 1604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1524952243
transform 1 0 1636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1524952243
transform 1 0 1556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1524952243
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1524952243
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1524952243
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1524952243
transform 1 0 1580 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1524952243
transform 1 0 1604 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1524952243
transform 1 0 1644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1524952243
transform 1 0 1716 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_551
timestamp 1524952243
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1524952243
transform 1 0 1692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1524952243
transform 1 0 1716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1524952243
transform 1 0 1684 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_531
timestamp 1524952243
transform 1 0 1692 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1524952243
transform 1 0 1764 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1524952243
transform 1 0 1852 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1524952243
transform 1 0 1756 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1524952243
transform 1 0 1796 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1524952243
transform 1 0 1756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1524952243
transform 1 0 1796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1524952243
transform 1 0 1852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1524952243
transform 1 0 1868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1524952243
transform 1 0 1740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1524952243
transform 1 0 1748 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1524952243
transform 1 0 1740 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_609
timestamp 1524952243
transform 1 0 1772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1524952243
transform 1 0 1860 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_467
timestamp 1524952243
transform 1 0 1908 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1524952243
transform 1 0 1908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1524952243
transform 1 0 1940 0 1 1405
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_10
timestamp 1524952243
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_10
timestamp 1524952243
transform 1 0 72 0 1 1370
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_37
timestamp 1524952243
transform -1 0 176 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_44
timestamp 1524952243
transform 1 0 176 0 1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_17
timestamp 1524952243
transform 1 0 192 0 1 1370
box -8 -3 34 105
use XOR2X1  XOR2X1_2
timestamp 1524952243
transform 1 0 224 0 1 1370
box -8 -3 64 105
use OAI21X1  OAI21X1_18
timestamp 1524952243
transform 1 0 280 0 1 1370
box -8 -3 34 105
use OR2X2  OR2X2_0
timestamp 1524952243
transform -1 0 344 0 1 1370
box -7 -3 35 105
use M3_M2  M3_M2_544
timestamp 1524952243
transform 1 0 364 0 1 1375
box -3 -3 3 3
use AND2X2  AND2X2_9
timestamp 1524952243
transform 1 0 344 0 1 1370
box -8 -3 40 105
use NAND2X1  NAND2X1_10
timestamp 1524952243
transform 1 0 376 0 1 1370
box -8 -3 32 105
use INVX2  INVX2_45
timestamp 1524952243
transform 1 0 400 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1524952243
transform 1 0 416 0 1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_1
timestamp 1524952243
transform 1 0 432 0 1 1370
box -8 -3 46 105
use BUFX2  BUFX2_3
timestamp 1524952243
transform -1 0 496 0 1 1370
box -5 -3 28 105
use OAI21X1  OAI21X1_19
timestamp 1524952243
transform 1 0 496 0 1 1370
box -8 -3 34 105
use M3_M2  M3_M2_545
timestamp 1524952243
transform 1 0 548 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_11
timestamp 1524952243
transform -1 0 552 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1524952243
transform 1 0 552 0 1 1370
box -8 -3 32 105
use M3_M2  M3_M2_546
timestamp 1524952243
transform 1 0 596 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1524952243
transform 1 0 660 0 1 1375
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_38
timestamp 1524952243
transform -1 0 672 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_548
timestamp 1524952243
transform 1 0 740 0 1 1375
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_39
timestamp 1524952243
transform 1 0 672 0 1 1370
box -8 -3 104 105
use NOR2X1  NOR2X1_9
timestamp 1524952243
transform 1 0 768 0 1 1370
box -8 -3 32 105
use M3_M2  M3_M2_549
timestamp 1524952243
transform 1 0 812 0 1 1375
box -3 -3 3 3
use OAI21X1  OAI21X1_26
timestamp 1524952243
transform 1 0 792 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1524952243
transform -1 0 856 0 1 1370
box -8 -3 34 105
use M3_M2  M3_M2_550
timestamp 1524952243
transform 1 0 940 0 1 1375
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_42
timestamp 1524952243
transform 1 0 856 0 1 1370
box -8 -3 104 105
use BUFX2  BUFX2_4
timestamp 1524952243
transform 1 0 952 0 1 1370
box -5 -3 28 105
use AOI22X1  AOI22X1_11
timestamp 1524952243
transform -1 0 1016 0 1 1370
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_43
timestamp 1524952243
transform 1 0 1016 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_53
timestamp 1524952243
transform -1 0 1128 0 1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_28
timestamp 1524952243
transform 1 0 1128 0 1 1370
box -8 -3 34 105
use XNOR2X1  XNOR2X1_0
timestamp 1524952243
transform 1 0 1160 0 1 1370
box -8 -3 64 105
use AND2X2  AND2X2_10
timestamp 1524952243
transform -1 0 1248 0 1 1370
box -8 -3 40 105
use M3_M2  M3_M2_551
timestamp 1524952243
transform 1 0 1308 0 1 1375
box -3 -3 3 3
use XOR2X1  XOR2X1_3
timestamp 1524952243
transform -1 0 1304 0 1 1370
box -8 -3 64 105
use AOI22X1  AOI22X1_12
timestamp 1524952243
transform 1 0 1304 0 1 1370
box -8 -3 46 105
use M3_M2  M3_M2_552
timestamp 1524952243
transform 1 0 1356 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_13
timestamp 1524952243
transform 1 0 1344 0 1 1370
box -8 -3 46 105
use AND2X2  AND2X2_11
timestamp 1524952243
transform -1 0 1416 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1524952243
transform 1 0 1416 0 1 1370
box -8 -3 40 105
use XNOR2X1  XNOR2X1_1
timestamp 1524952243
transform -1 0 1504 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1524952243
transform 1 0 1504 0 1 1370
box -8 -3 64 105
use AOI22X1  AOI22X1_14
timestamp 1524952243
transform 1 0 1560 0 1 1370
box -8 -3 46 105
use XNOR2X1  XNOR2X1_2
timestamp 1524952243
transform 1 0 1600 0 1 1370
box -8 -3 64 105
use AND2X2  AND2X2_13
timestamp 1524952243
transform -1 0 1688 0 1 1370
box -8 -3 40 105
use XOR2X1  XOR2X1_5
timestamp 1524952243
transform 1 0 1688 0 1 1370
box -8 -3 64 105
use INVX2  INVX2_54
timestamp 1524952243
transform 1 0 1744 0 1 1370
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_44
timestamp 1524952243
transform 1 0 1760 0 1 1370
box -8 -3 104 105
use AND2X2  AND2X2_14
timestamp 1524952243
transform 1 0 1856 0 1 1370
box -8 -3 40 105
use XNOR2X1  XNOR2X1_3
timestamp 1524952243
transform -1 0 1944 0 1 1370
box -8 -3 64 105
use top_module_VIA0  top_module_VIA0_11
timestamp 1524952243
transform 1 0 1970 0 1 1370
box -10 -3 10 3
use M3_M2  M3_M2_553
timestamp 1524952243
transform 1 0 116 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_617
timestamp 1524952243
transform 1 0 76 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1524952243
transform 1 0 100 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_565
timestamp 1524952243
transform 1 0 124 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_619
timestamp 1524952243
transform 1 0 124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1524952243
transform 1 0 132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1524952243
transform 1 0 148 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_616
timestamp 1524952243
transform 1 0 92 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1524952243
transform 1 0 108 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_679
timestamp 1524952243
transform 1 0 116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1524952243
transform 1 0 124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1524952243
transform 1 0 148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1524952243
transform 1 0 92 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_673
timestamp 1524952243
transform 1 0 68 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_613
timestamp 1524952243
transform 1 0 164 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_579
timestamp 1524952243
transform 1 0 172 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1524952243
transform 1 0 204 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1524952243
transform 1 0 204 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_622
timestamp 1524952243
transform 1 0 188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1524952243
transform 1 0 196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1524952243
transform 1 0 204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1524952243
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_618
timestamp 1524952243
transform 1 0 180 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1524952243
transform 1 0 228 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_683
timestamp 1524952243
transform 1 0 204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1524952243
transform 1 0 212 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_642
timestamp 1524952243
transform 1 0 164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1524952243
transform 1 0 188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1524952243
transform 1 0 172 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1524952243
transform 1 0 180 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_748
timestamp 1524952243
transform 1 0 228 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1524952243
transform 1 0 228 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_685
timestamp 1524952243
transform 1 0 244 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_619
timestamp 1524952243
transform 1 0 252 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1524952243
transform 1 0 284 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_625
timestamp 1524952243
transform 1 0 284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1524952243
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1524952243
transform 1 0 252 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_620
timestamp 1524952243
transform 1 0 276 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_687
timestamp 1524952243
transform 1 0 284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1524952243
transform 1 0 276 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_644
timestamp 1524952243
transform 1 0 284 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_770
timestamp 1524952243
transform 1 0 268 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_675
timestamp 1524952243
transform 1 0 252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1524952243
transform 1 0 268 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1524952243
transform 1 0 212 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1524952243
transform 1 0 236 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1524952243
transform 1 0 276 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1524952243
transform 1 0 300 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1524952243
transform 1 0 292 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1524952243
transform 1 0 292 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1524952243
transform 1 0 300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1524952243
transform 1 0 308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1524952243
transform 1 0 324 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_622
timestamp 1524952243
transform 1 0 332 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_626
timestamp 1524952243
transform 1 0 428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1524952243
transform 1 0 348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1524952243
transform 1 0 324 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_645
timestamp 1524952243
transform 1 0 332 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1524952243
transform 1 0 356 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_692
timestamp 1524952243
transform 1 0 396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1524952243
transform 1 0 444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1524952243
transform 1 0 340 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1524952243
transform 1 0 308 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_771
timestamp 1524952243
transform 1 0 316 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1524952243
transform 1 0 324 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1524952243
transform 1 0 412 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1524952243
transform 1 0 428 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1524952243
transform 1 0 364 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1524952243
transform 1 0 388 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1524952243
transform 1 0 428 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1524952243
transform 1 0 572 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1524952243
transform 1 0 476 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1524952243
transform 1 0 556 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1524952243
transform 1 0 564 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_627
timestamp 1524952243
transform 1 0 548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1524952243
transform 1 0 564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1524952243
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1524952243
transform 1 0 468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1524952243
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_624
timestamp 1524952243
transform 1 0 548 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_753
timestamp 1524952243
transform 1 0 460 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1524952243
transform 1 0 460 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1524952243
transform 1 0 596 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_629
timestamp 1524952243
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1524952243
transform 1 0 572 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_648
timestamp 1524952243
transform 1 0 564 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1524952243
transform 1 0 540 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1524952243
transform 1 0 580 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1524952243
transform 1 0 604 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_630
timestamp 1524952243
transform 1 0 604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1524952243
transform 1 0 612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1524952243
transform 1 0 596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1524952243
transform 1 0 580 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1524952243
transform 1 0 572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1524952243
transform 1 0 580 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_614
timestamp 1524952243
transform 1 0 644 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_585
timestamp 1524952243
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1524952243
transform 1 0 684 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_632
timestamp 1524952243
transform 1 0 636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1524952243
transform 1 0 652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1524952243
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_649
timestamp 1524952243
transform 1 0 612 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1524952243
transform 1 0 636 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1524952243
transform 1 0 636 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_681
timestamp 1524952243
transform 1 0 620 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1524952243
transform 1 0 660 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_634
timestamp 1524952243
transform 1 0 668 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1524952243
transform 1 0 684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1524952243
transform 1 0 660 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_627
timestamp 1524952243
transform 1 0 676 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_615
timestamp 1524952243
transform 1 0 716 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1524952243
transform 1 0 724 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1524952243
transform 1 0 708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1524952243
transform 1 0 684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1524952243
transform 1 0 692 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_650
timestamp 1524952243
transform 1 0 660 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1524952243
transform 1 0 684 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1524952243
transform 1 0 708 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_756
timestamp 1524952243
transform 1 0 708 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1524952243
transform 1 0 748 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_616
timestamp 1524952243
transform 1 0 772 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1524952243
transform 1 0 748 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1524952243
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_605
timestamp 1524952243
transform 1 0 772 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_703
timestamp 1524952243
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1524952243
transform 1 0 748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_652
timestamp 1524952243
transform 1 0 732 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1524952243
transform 1 0 692 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1524952243
transform 1 0 716 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1524952243
transform 1 0 732 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1524952243
transform 1 0 668 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1524952243
transform 1 0 716 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1524952243
transform 1 0 764 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1524952243
transform 1 0 764 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_556
timestamp 1524952243
transform 1 0 828 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1524952243
transform 1 0 812 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1524952243
transform 1 0 804 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1524952243
transform 1 0 836 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1524952243
transform 1 0 948 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1524952243
transform 1 0 964 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1524952243
transform 1 0 940 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1524952243
transform 1 0 1084 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1524952243
transform 1 0 1068 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1524952243
transform 1 0 1020 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_638
timestamp 1524952243
transform 1 0 820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1524952243
transform 1 0 828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1524952243
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1524952243
transform 1 0 940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1524952243
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1524952243
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1524952243
transform 1 0 980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1524952243
transform 1 0 988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1524952243
transform 1 0 788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1524952243
transform 1 0 804 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1524952243
transform 1 0 788 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1524952243
transform 1 0 820 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1524952243
transform 1 0 828 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_631
timestamp 1524952243
transform 1 0 852 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_708
timestamp 1524952243
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1524952243
transform 1 0 916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1524952243
transform 1 0 820 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1524952243
transform 1 0 828 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1524952243
transform 1 0 852 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1524952243
transform 1 0 852 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1524952243
transform 1 0 828 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_710
timestamp 1524952243
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_632
timestamp 1524952243
transform 1 0 980 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1524952243
transform 1 0 1116 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1524952243
transform 1 0 1132 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1524952243
transform 1 0 1148 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_646
timestamp 1524952243
transform 1 0 1020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1524952243
transform 1 0 1108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1524952243
transform 1 0 988 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1524952243
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1524952243
transform 1 0 1044 0 1 1324
box -2 -2 2 2
use M3_M2  M3_M2_633
timestamp 1524952243
transform 1 0 1092 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1524952243
transform 1 0 1132 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1524952243
transform 1 0 1188 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1524952243
transform 1 0 1156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1524952243
transform 1 0 1172 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_648
timestamp 1524952243
transform 1 0 1140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1524952243
transform 1 0 1148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1524952243
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1524952243
transform 1 0 1108 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1524952243
transform 1 0 1004 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1524952243
transform 1 0 1044 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_715
timestamp 1524952243
transform 1 0 1132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1524952243
transform 1 0 1124 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_634
timestamp 1524952243
transform 1 0 1140 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_716
timestamp 1524952243
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_562
timestamp 1524952243
transform 1 0 1252 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1524952243
transform 1 0 1204 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1524952243
transform 1 0 1244 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1524952243
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1524952243
transform 1 0 1196 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1524952243
transform 1 0 1268 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_651
timestamp 1524952243
transform 1 0 1268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1524952243
transform 1 0 1196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1524952243
transform 1 0 1212 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_635
timestamp 1524952243
transform 1 0 1236 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_719
timestamp 1524952243
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1524952243
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1524952243
transform 1 0 1204 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1524952243
transform 1 0 1188 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1524952243
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_577
timestamp 1524952243
transform 1 0 1356 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1524952243
transform 1 0 1348 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1524952243
transform 1 0 1348 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_653
timestamp 1524952243
transform 1 0 1356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1524952243
transform 1 0 1364 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_610
timestamp 1524952243
transform 1 0 1372 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_655
timestamp 1524952243
transform 1 0 1388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1524952243
transform 1 0 1396 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_595
timestamp 1524952243
transform 1 0 1452 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_657
timestamp 1524952243
transform 1 0 1444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1524952243
transform 1 0 1452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1524952243
transform 1 0 1316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1524952243
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1524952243
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1524952243
transform 1 0 1356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1524952243
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1524952243
transform 1 0 1388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1524952243
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1524952243
transform 1 0 1316 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1524952243
transform 1 0 1292 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1524952243
transform 1 0 1324 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1524952243
transform 1 0 1388 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1524952243
transform 1 0 1412 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1524952243
transform 1 0 1364 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1524952243
transform 1 0 1388 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1524952243
transform 1 0 1580 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1524952243
transform 1 0 1596 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1524952243
transform 1 0 1572 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1524952243
transform 1 0 1484 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1524952243
transform 1 0 1516 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1524952243
transform 1 0 1548 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_659
timestamp 1524952243
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1524952243
transform 1 0 1484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1524952243
transform 1 0 1508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1524952243
transform 1 0 1516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1524952243
transform 1 0 1524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1524952243
transform 1 0 1460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1524952243
transform 1 0 1476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1524952243
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1524952243
transform 1 0 1476 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_611
timestamp 1524952243
transform 1 0 1532 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_664
timestamp 1524952243
transform 1 0 1540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1524952243
transform 1 0 1548 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_612
timestamp 1524952243
transform 1 0 1556 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_666
timestamp 1524952243
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1524952243
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1524952243
transform 1 0 1588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1524952243
transform 1 0 1596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1524952243
transform 1 0 1516 0 1 1324
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1524952243
transform 1 0 1532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1524952243
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1524952243
transform 1 0 1556 0 1 1324
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1524952243
transform 1 0 1572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1524952243
transform 1 0 1596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1524952243
transform 1 0 1508 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1524952243
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_613
timestamp 1524952243
transform 1 0 1636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1524952243
transform 1 0 1668 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_671
timestamp 1524952243
transform 1 0 1644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1524952243
transform 1 0 1668 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1524952243
transform 1 0 1612 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_735
timestamp 1524952243
transform 1 0 1620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_658
timestamp 1524952243
transform 1 0 1556 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1524952243
transform 1 0 1596 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_764
timestamp 1524952243
transform 1 0 1612 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_698
timestamp 1524952243
transform 1 0 1540 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1524952243
transform 1 0 1588 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1524952243
transform 1 0 1564 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1524952243
transform 1 0 1580 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1524952243
transform 1 0 1628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1524952243
transform 1 0 1740 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1524952243
transform 1 0 1740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1524952243
transform 1 0 1684 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_637
timestamp 1524952243
transform 1 0 1708 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_674
timestamp 1524952243
transform 1 0 1796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1524952243
transform 1 0 1716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1524952243
transform 1 0 1732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1524952243
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1524952243
transform 1 0 1788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1524952243
transform 1 0 1644 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1524952243
transform 1 0 1652 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1524952243
transform 1 0 1676 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1524952243
transform 1 0 1668 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_638
timestamp 1524952243
transform 1 0 1796 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1524952243
transform 1 0 1884 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_675
timestamp 1524952243
transform 1 0 1844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1524952243
transform 1 0 1820 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_614
timestamp 1524952243
transform 1 0 1860 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_676
timestamp 1524952243
transform 1 0 1884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1524952243
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_639
timestamp 1524952243
transform 1 0 1868 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_768
timestamp 1524952243
transform 1 0 1852 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_687
timestamp 1524952243
transform 1 0 1820 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1524952243
transform 1 0 1860 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1524952243
transform 1 0 1868 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_615
timestamp 1524952243
transform 1 0 1892 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_677
timestamp 1524952243
transform 1 0 1916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1524952243
transform 1 0 1940 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_640
timestamp 1524952243
transform 1 0 1916 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_743
timestamp 1524952243
transform 1 0 1924 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_641
timestamp 1524952243
transform 1 0 1948 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_769
timestamp 1524952243
transform 1 0 1940 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1524952243
transform 1 0 1940 0 1 1305
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_12
timestamp 1524952243
transform 1 0 24 0 1 1270
box -10 -3 10 3
use NAND2X1  NAND2X1_13
timestamp 1524952243
transform 1 0 72 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_20
timestamp 1524952243
transform -1 0 128 0 -1 1370
box -8 -3 34 105
use INVX2  INVX2_47
timestamp 1524952243
transform 1 0 128 0 -1 1370
box -9 -3 26 105
use NOR2X1  NOR2X1_10
timestamp 1524952243
transform -1 0 168 0 -1 1370
box -8 -3 32 105
use AOI21X1  AOI21X1_6
timestamp 1524952243
transform -1 0 200 0 -1 1370
box -7 -3 39 105
use OAI21X1  OAI21X1_21
timestamp 1524952243
transform 1 0 200 0 -1 1370
box -8 -3 34 105
use INVX2  INVX2_48
timestamp 1524952243
transform 1 0 232 0 -1 1370
box -9 -3 26 105
use NAND3X1  NAND3X1_10
timestamp 1524952243
transform 1 0 248 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_49
timestamp 1524952243
transform 1 0 280 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1524952243
transform 1 0 296 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_700
timestamp 1524952243
transform 1 0 348 0 1 1275
box -3 -3 3 3
use NAND3X1  NAND3X1_11
timestamp 1524952243
transform 1 0 312 0 -1 1370
box -8 -3 40 105
use M3_M2  M3_M2_701
timestamp 1524952243
transform 1 0 364 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1524952243
transform 1 0 380 0 1 1275
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_40
timestamp 1524952243
transform -1 0 440 0 -1 1370
box -8 -3 104 105
use NAND2X1  NAND2X1_14
timestamp 1524952243
transform 1 0 440 0 -1 1370
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_41
timestamp 1524952243
transform -1 0 560 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_51
timestamp 1524952243
transform 1 0 560 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_703
timestamp 1524952243
transform 1 0 596 0 1 1275
box -3 -3 3 3
use OAI21X1  OAI21X1_22
timestamp 1524952243
transform -1 0 608 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1524952243
transform 1 0 608 0 -1 1370
box -8 -3 34 105
use NOR2X1  NOR2X1_11
timestamp 1524952243
transform 1 0 640 0 -1 1370
box -8 -3 32 105
use INVX2  INVX2_52
timestamp 1524952243
transform 1 0 664 0 -1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_24
timestamp 1524952243
transform 1 0 680 0 -1 1370
box -8 -3 34 105
use NOR2X1  NOR2X1_12
timestamp 1524952243
transform 1 0 712 0 -1 1370
box -8 -3 32 105
use M3_M2  M3_M2_704
timestamp 1524952243
transform 1 0 764 0 1 1275
box -3 -3 3 3
use OAI21X1  OAI21X1_25
timestamp 1524952243
transform 1 0 736 0 -1 1370
box -8 -3 34 105
use NOR2X1  NOR2X1_13
timestamp 1524952243
transform 1 0 768 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_29
timestamp 1524952243
transform 1 0 792 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1524952243
transform 1 0 824 0 -1 1370
box -8 -3 34 105
use M3_M2  M3_M2_705
timestamp 1524952243
transform 1 0 900 0 1 1275
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_45
timestamp 1524952243
transform -1 0 952 0 -1 1370
box -8 -3 104 105
use AOI22X1  AOI22X1_15
timestamp 1524952243
transform -1 0 992 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_55
timestamp 1524952243
transform 1 0 992 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_706
timestamp 1524952243
transform 1 0 1108 0 1 1275
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_46
timestamp 1524952243
transform 1 0 1008 0 -1 1370
box -8 -3 104 105
use M3_M2  M3_M2_707
timestamp 1524952243
transform 1 0 1132 0 1 1275
box -3 -3 3 3
use INVX2  INVX2_56
timestamp 1524952243
transform 1 0 1104 0 -1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_15
timestamp 1524952243
transform -1 0 1144 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_31
timestamp 1524952243
transform 1 0 1144 0 -1 1370
box -8 -3 34 105
use M3_M2  M3_M2_708
timestamp 1524952243
transform 1 0 1204 0 1 1275
box -3 -3 3 3
use NAND3X1  NAND3X1_12
timestamp 1524952243
transform -1 0 1208 0 -1 1370
box -8 -3 40 105
use XNOR2X1  XNOR2X1_4
timestamp 1524952243
transform 1 0 1208 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1524952243
transform 1 0 1264 0 -1 1370
box -8 -3 64 105
use M3_M2  M3_M2_709
timestamp 1524952243
transform 1 0 1348 0 1 1275
box -3 -3 3 3
use AND2X2  AND2X2_15
timestamp 1524952243
transform -1 0 1352 0 -1 1370
box -8 -3 40 105
use AOI22X1  AOI22X1_16
timestamp 1524952243
transform 1 0 1352 0 -1 1370
box -8 -3 46 105
use XOR2X1  XOR2X1_7
timestamp 1524952243
transform -1 0 1448 0 -1 1370
box -8 -3 64 105
use OAI21X1  OAI21X1_32
timestamp 1524952243
transform 1 0 1448 0 -1 1370
box -8 -3 34 105
use M3_M2  M3_M2_710
timestamp 1524952243
transform 1 0 1524 0 1 1275
box -3 -3 3 3
use OAI21X1  OAI21X1_33
timestamp 1524952243
transform 1 0 1480 0 -1 1370
box -8 -3 34 105
use AOI22X1  AOI22X1_17
timestamp 1524952243
transform 1 0 1512 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1524952243
transform 1 0 1552 0 -1 1370
box -8 -3 46 105
use NAND2X1  NAND2X1_16
timestamp 1524952243
transform 1 0 1592 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_34
timestamp 1524952243
transform 1 0 1616 0 -1 1370
box -8 -3 34 105
use NAND3X1  NAND3X1_13
timestamp 1524952243
transform -1 0 1680 0 -1 1370
box -8 -3 40 105
use XNOR2X1  XNOR2X1_5
timestamp 1524952243
transform 1 0 1680 0 -1 1370
box -8 -3 64 105
use M3_M2  M3_M2_711
timestamp 1524952243
transform 1 0 1764 0 1 1275
box -3 -3 3 3
use XOR2X1  XOR2X1_8
timestamp 1524952243
transform 1 0 1736 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1524952243
transform 1 0 1792 0 -1 1370
box -8 -3 64 105
use NAND3X1  NAND3X1_14
timestamp 1524952243
transform 1 0 1848 0 -1 1370
box -8 -3 40 105
use OAI21X1  OAI21X1_35
timestamp 1524952243
transform -1 0 1912 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1524952243
transform 1 0 1912 0 -1 1370
box -8 -3 34 105
use top_module_VIA0  top_module_VIA0_13
timestamp 1524952243
transform 1 0 1994 0 1 1270
box -10 -3 10 3
use M3_M2  M3_M2_712
timestamp 1524952243
transform 1 0 164 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1524952243
transform 1 0 124 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1524952243
transform 1 0 68 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1524952243
transform 1 0 132 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_775
timestamp 1524952243
transform 1 0 196 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1524952243
transform 1 0 172 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1524952243
transform 1 0 188 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1524952243
transform 1 0 68 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1524952243
transform 1 0 116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1524952243
transform 1 0 156 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_837
timestamp 1524952243
transform 1 0 84 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1524952243
transform 1 0 116 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1524952243
transform 1 0 156 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_790
timestamp 1524952243
transform 1 0 188 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1524952243
transform 1 0 196 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_856
timestamp 1524952243
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1524952243
transform 1 0 204 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1524952243
transform 1 0 220 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1524952243
transform 1 0 220 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1524952243
transform 1 0 228 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_913
timestamp 1524952243
transform 1 0 228 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1524952243
transform 1 0 228 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1524952243
transform 1 0 252 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1524952243
transform 1 0 244 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_792
timestamp 1524952243
transform 1 0 252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1524952243
transform 1 0 244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1524952243
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_759
timestamp 1524952243
transform 1 0 268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1524952243
transform 1 0 292 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1524952243
transform 1 0 308 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1524952243
transform 1 0 300 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1524952243
transform 1 0 292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1524952243
transform 1 0 300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1524952243
transform 1 0 284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1524952243
transform 1 0 268 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1524952243
transform 1 0 276 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_841
timestamp 1524952243
transform 1 0 276 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1524952243
transform 1 0 340 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1524952243
transform 1 0 332 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_779
timestamp 1524952243
transform 1 0 348 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_762
timestamp 1524952243
transform 1 0 356 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1524952243
transform 1 0 316 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_795
timestamp 1524952243
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1524952243
transform 1 0 308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1524952243
transform 1 0 316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1524952243
transform 1 0 316 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_786
timestamp 1524952243
transform 1 0 348 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_796
timestamp 1524952243
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1524952243
transform 1 0 348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_842
timestamp 1524952243
transform 1 0 340 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1524952243
transform 1 0 388 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1524952243
transform 1 0 420 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1524952243
transform 1 0 380 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1524952243
transform 1 0 404 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1524952243
transform 1 0 380 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1524952243
transform 1 0 404 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1524952243
transform 1 0 388 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_797
timestamp 1524952243
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1524952243
transform 1 0 404 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1524952243
transform 1 0 428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1524952243
transform 1 0 364 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1524952243
transform 1 0 380 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_864
timestamp 1524952243
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_809
timestamp 1524952243
transform 1 0 404 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1524952243
transform 1 0 452 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_865
timestamp 1524952243
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1524952243
transform 1 0 436 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_821
timestamp 1524952243
transform 1 0 380 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1524952243
transform 1 0 372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1524952243
transform 1 0 444 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1524952243
transform 1 0 468 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1524952243
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1524952243
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1524952243
transform 1 0 444 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1524952243
transform 1 0 452 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_844
timestamp 1524952243
transform 1 0 436 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1524952243
transform 1 0 460 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1524952243
transform 1 0 500 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1524952243
transform 1 0 484 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1524952243
transform 1 0 500 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_781
timestamp 1524952243
transform 1 0 508 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1524952243
transform 1 0 484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1524952243
transform 1 0 492 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_811
timestamp 1524952243
transform 1 0 492 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1524952243
transform 1 0 476 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1524952243
transform 1 0 556 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1524952243
transform 1 0 548 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1524952243
transform 1 0 532 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_782
timestamp 1524952243
transform 1 0 548 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1524952243
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_787
timestamp 1524952243
transform 1 0 516 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1524952243
transform 1 0 564 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_802
timestamp 1524952243
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1524952243
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1524952243
transform 1 0 548 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_788
timestamp 1524952243
transform 1 0 564 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_869
timestamp 1524952243
transform 1 0 524 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_812
timestamp 1524952243
transform 1 0 548 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1524952243
transform 1 0 532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1524952243
transform 1 0 548 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1524952243
transform 1 0 604 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_805
timestamp 1524952243
transform 1 0 596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1524952243
transform 1 0 620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1524952243
transform 1 0 580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1524952243
transform 1 0 588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1524952243
transform 1 0 604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1524952243
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_823
timestamp 1524952243
transform 1 0 620 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1524952243
transform 1 0 644 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1524952243
transform 1 0 660 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1524952243
transform 1 0 636 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1524952243
transform 1 0 636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1524952243
transform 1 0 636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1524952243
transform 1 0 660 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1524952243
transform 1 0 724 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1524952243
transform 1 0 652 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1524952243
transform 1 0 692 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1524952243
transform 1 0 708 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_808
timestamp 1524952243
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1524952243
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_789
timestamp 1524952243
transform 1 0 684 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_810
timestamp 1524952243
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1524952243
transform 1 0 732 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_824
timestamp 1524952243
transform 1 0 708 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1524952243
transform 1 0 756 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_811
timestamp 1524952243
transform 1 0 780 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_791
timestamp 1524952243
transform 1 0 804 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1524952243
transform 1 0 828 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_812
timestamp 1524952243
transform 1 0 836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1524952243
transform 1 0 844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1524952243
transform 1 0 756 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_813
timestamp 1524952243
transform 1 0 820 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1524952243
transform 1 0 756 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1524952243
transform 1 0 836 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1524952243
transform 1 0 748 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1524952243
transform 1 0 780 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1524952243
transform 1 0 804 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_814
timestamp 1524952243
transform 1 0 852 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_793
timestamp 1524952243
transform 1 0 860 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_877
timestamp 1524952243
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_726
timestamp 1524952243
transform 1 0 876 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1524952243
transform 1 0 876 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1524952243
transform 1 0 908 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1524952243
transform 1 0 924 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1524952243
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1524952243
transform 1 0 876 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_794
timestamp 1524952243
transform 1 0 884 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1524952243
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1524952243
transform 1 0 908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1524952243
transform 1 0 916 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1524952243
transform 1 0 988 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1524952243
transform 1 0 956 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_820
timestamp 1524952243
transform 1 0 932 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_795
timestamp 1524952243
transform 1 0 948 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_821
timestamp 1524952243
transform 1 0 956 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_796
timestamp 1524952243
transform 1 0 964 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_822
timestamp 1524952243
transform 1 0 972 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_797
timestamp 1524952243
transform 1 0 980 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1524952243
transform 1 0 1100 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1524952243
transform 1 0 1004 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1524952243
transform 1 0 1044 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_823
timestamp 1524952243
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1524952243
transform 1 0 1004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1524952243
transform 1 0 1044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1524952243
transform 1 0 884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1524952243
transform 1 0 900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1524952243
transform 1 0 908 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_814
timestamp 1524952243
transform 1 0 916 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1524952243
transform 1 0 932 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1524952243
transform 1 0 884 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_881
timestamp 1524952243
transform 1 0 964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1524952243
transform 1 0 980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1524952243
transform 1 0 988 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_827
timestamp 1524952243
transform 1 0 964 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1524952243
transform 1 0 1092 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_826
timestamp 1524952243
transform 1 0 1100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1524952243
transform 1 0 1108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1524952243
transform 1 0 1020 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_828
timestamp 1524952243
transform 1 0 1036 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1524952243
transform 1 0 1124 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1524952243
transform 1 0 1124 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_828
timestamp 1524952243
transform 1 0 1116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1524952243
transform 1 0 1124 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1524952243
transform 1 0 1148 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1524952243
transform 1 0 1140 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_830
timestamp 1524952243
transform 1 0 1140 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1524952243
transform 1 0 1164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1524952243
transform 1 0 1180 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_831
timestamp 1524952243
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1524952243
transform 1 0 1156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1524952243
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1524952243
transform 1 0 1180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1524952243
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_816
timestamp 1524952243
transform 1 0 1148 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1524952243
transform 1 0 1188 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_886
timestamp 1524952243
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1524952243
transform 1 0 1188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1524952243
transform 1 0 1196 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_829
timestamp 1524952243
transform 1 0 1172 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1524952243
transform 1 0 1260 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_835
timestamp 1524952243
transform 1 0 1204 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_800
timestamp 1524952243
transform 1 0 1236 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_836
timestamp 1524952243
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1524952243
transform 1 0 1284 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1524952243
transform 1 0 1300 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_817
timestamp 1524952243
transform 1 0 1204 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_889
timestamp 1524952243
transform 1 0 1220 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_818
timestamp 1524952243
transform 1 0 1308 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1524952243
transform 1 0 1324 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1524952243
transform 1 0 1372 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1524952243
transform 1 0 1332 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1524952243
transform 1 0 1404 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1524952243
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1524952243
transform 1 0 1332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1524952243
transform 1 0 1348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1524952243
transform 1 0 1316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1524952243
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_830
timestamp 1524952243
transform 1 0 1244 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1524952243
transform 1 0 1308 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_852
timestamp 1524952243
transform 1 0 1300 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1524952243
transform 1 0 1332 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1524952243
transform 1 0 1380 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_783
timestamp 1524952243
transform 1 0 1412 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1524952243
transform 1 0 1388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1524952243
transform 1 0 1404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1524952243
transform 1 0 1380 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_853
timestamp 1524952243
transform 1 0 1340 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_776
timestamp 1524952243
transform 1 0 1436 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_778
timestamp 1524952243
transform 1 0 1428 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_893
timestamp 1524952243
transform 1 0 1428 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_750
timestamp 1524952243
transform 1 0 1460 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_784
timestamp 1524952243
transform 1 0 1460 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1524952243
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1524952243
transform 1 0 1468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1524952243
transform 1 0 1468 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_832
timestamp 1524952243
transform 1 0 1444 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_785
timestamp 1524952243
transform 1 0 1484 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1524952243
transform 1 0 1516 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1524952243
transform 1 0 1508 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1524952243
transform 1 0 1540 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1524952243
transform 1 0 1532 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_845
timestamp 1524952243
transform 1 0 1532 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1524952243
transform 1 0 1540 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_895
timestamp 1524952243
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_819
timestamp 1524952243
transform 1 0 1532 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1524952243
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1524952243
transform 1 0 1620 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1524952243
transform 1 0 1588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1524952243
transform 1 0 1612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1524952243
transform 1 0 1548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1524952243
transform 1 0 1508 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_833
timestamp 1524952243
transform 1 0 1516 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1524952243
transform 1 0 1508 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1524952243
transform 1 0 1556 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_897
timestamp 1524952243
transform 1 0 1564 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_834
timestamp 1524952243
transform 1 0 1548 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_921
timestamp 1524952243
transform 1 0 1556 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1524952243
transform 1 0 1564 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_898
timestamp 1524952243
transform 1 0 1612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1524952243
transform 1 0 1620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1524952243
transform 1 0 1612 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_786
timestamp 1524952243
transform 1 0 1644 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1524952243
transform 1 0 1676 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_848
timestamp 1524952243
transform 1 0 1668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1524952243
transform 1 0 1700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1524952243
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1524952243
transform 1 0 1652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1524952243
transform 1 0 1700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1524952243
transform 1 0 1708 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_836
timestamp 1524952243
transform 1 0 1644 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1524952243
transform 1 0 1708 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1524952243
transform 1 0 1748 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1524952243
transform 1 0 1788 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_850
timestamp 1524952243
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1524952243
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1524952243
transform 1 0 1732 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1524952243
transform 1 0 1724 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_783
timestamp 1524952243
transform 1 0 1812 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_905
timestamp 1524952243
transform 1 0 1780 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1524952243
transform 1 0 1796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1524952243
transform 1 0 1812 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1524952243
transform 1 0 1724 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1524952243
transform 1 0 1772 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_923
timestamp 1524952243
transform 1 0 1804 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_859
timestamp 1524952243
transform 1 0 1804 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1524952243
transform 1 0 1884 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1524952243
transform 1 0 1924 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1524952243
transform 1 0 1868 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1524952243
transform 1 0 1924 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1524952243
transform 1 0 1884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1524952243
transform 1 0 1892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1524952243
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1524952243
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1524952243
transform 1 0 1924 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_854
timestamp 1524952243
transform 1 0 1940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1524952243
transform 1 0 1916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1524952243
transform 1 0 1948 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1524952243
transform 1 0 1860 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1524952243
transform 1 0 1892 0 1 1185
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_14
timestamp 1524952243
transform 1 0 48 0 1 1170
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_47
timestamp 1524952243
transform -1 0 168 0 1 1170
box -8 -3 104 105
use NAND3X1  NAND3X1_15
timestamp 1524952243
transform -1 0 200 0 1 1170
box -8 -3 40 105
use M3_M2  M3_M2_862
timestamp 1524952243
transform 1 0 220 0 1 1175
box -3 -3 3 3
use NOR2X1  NOR2X1_14
timestamp 1524952243
transform 1 0 200 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1524952243
transform 1 0 224 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1524952243
transform -1 0 272 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_863
timestamp 1524952243
transform 1 0 284 0 1 1175
box -3 -3 3 3
use NOR2X1  NOR2X1_17
timestamp 1524952243
transform 1 0 272 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1524952243
transform -1 0 320 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_37
timestamp 1524952243
transform 1 0 320 0 1 1170
box -8 -3 34 105
use INVX2  INVX2_57
timestamp 1524952243
transform -1 0 368 0 1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_38
timestamp 1524952243
transform 1 0 368 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_864
timestamp 1524952243
transform 1 0 420 0 1 1175
box -3 -3 3 3
use NAND2X1  NAND2X1_17
timestamp 1524952243
transform -1 0 424 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1524952243
transform -1 0 448 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_865
timestamp 1524952243
transform 1 0 460 0 1 1175
box -3 -3 3 3
use NOR2X1  NOR2X1_20
timestamp 1524952243
transform 1 0 448 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_866
timestamp 1524952243
transform 1 0 484 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_58
timestamp 1524952243
transform 1 0 472 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1524952243
transform -1 0 504 0 1 1170
box -9 -3 26 105
use NAND2X1  NAND2X1_18
timestamp 1524952243
transform -1 0 528 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1524952243
transform 1 0 528 0 1 1170
box -8 -3 32 105
use BUFX2  BUFX2_5
timestamp 1524952243
transform 1 0 552 0 1 1170
box -5 -3 28 105
use AOI22X1  AOI22X1_19
timestamp 1524952243
transform -1 0 616 0 1 1170
box -8 -3 46 105
use INVX2  INVX2_60
timestamp 1524952243
transform 1 0 616 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1524952243
transform 1 0 632 0 1 1170
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_49
timestamp 1524952243
transform -1 0 744 0 1 1170
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_50
timestamp 1524952243
transform 1 0 744 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_62
timestamp 1524952243
transform 1 0 840 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1524952243
transform 1 0 856 0 1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_20
timestamp 1524952243
transform 1 0 872 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_867
timestamp 1524952243
transform 1 0 940 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_64
timestamp 1524952243
transform 1 0 912 0 1 1170
box -9 -3 26 105
use BUFX2  BUFX2_6
timestamp 1524952243
transform 1 0 928 0 1 1170
box -5 -3 28 105
use AOI22X1  AOI22X1_21
timestamp 1524952243
transform -1 0 992 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_868
timestamp 1524952243
transform 1 0 1012 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1524952243
transform 1 0 1052 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_65
timestamp 1524952243
transform 1 0 992 0 1 1170
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_51
timestamp 1524952243
transform 1 0 1008 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_870
timestamp 1524952243
transform 1 0 1116 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_66
timestamp 1524952243
transform 1 0 1104 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1524952243
transform 1 0 1120 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1524952243
transform 1 0 1136 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_871
timestamp 1524952243
transform 1 0 1180 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_2
timestamp 1524952243
transform 1 0 1152 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_872
timestamp 1524952243
transform 1 0 1204 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_69
timestamp 1524952243
transform 1 0 1192 0 1 1170
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_52
timestamp 1524952243
transform 1 0 1208 0 1 1170
box -8 -3 104 105
use NOR2X1  NOR2X1_21
timestamp 1524952243
transform 1 0 1304 0 1 1170
box -8 -3 32 105
use XNOR2X1  XNOR2X1_6
timestamp 1524952243
transform -1 0 1384 0 1 1170
box -8 -3 64 105
use AND2X2  AND2X2_16
timestamp 1524952243
transform -1 0 1416 0 1 1170
box -8 -3 40 105
use FILL  FILL_11
timestamp 1524952243
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_12
timestamp 1524952243
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1524952243
transform 1 0 1432 0 1 1170
box -8 -3 40 105
use NAND2X1  NAND2X1_20
timestamp 1524952243
transform 1 0 1464 0 1 1170
box -8 -3 32 105
use INVX2  INVX2_70
timestamp 1524952243
transform -1 0 1504 0 1 1170
box -9 -3 26 105
use AOI21X1  AOI21X1_7
timestamp 1524952243
transform -1 0 1536 0 1 1170
box -7 -3 39 105
use NOR2X1  NOR2X1_22
timestamp 1524952243
transform -1 0 1560 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_873
timestamp 1524952243
transform 1 0 1604 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_10
timestamp 1524952243
transform 1 0 1560 0 1 1170
box -8 -3 64 105
use OAI21X1  OAI21X1_39
timestamp 1524952243
transform 1 0 1616 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_874
timestamp 1524952243
transform 1 0 1700 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_11
timestamp 1524952243
transform -1 0 1704 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_875
timestamp 1524952243
transform 1 0 1732 0 1 1175
box -3 -3 3 3
use NOR2X1  NOR2X1_23
timestamp 1524952243
transform -1 0 1728 0 1 1170
box -8 -3 32 105
use XOR2X1  XOR2X1_12
timestamp 1524952243
transform -1 0 1784 0 1 1170
box -8 -3 64 105
use NOR2X1  NOR2X1_24
timestamp 1524952243
transform -1 0 1808 0 1 1170
box -8 -3 32 105
use XNOR2X1  XNOR2X1_7
timestamp 1524952243
transform 1 0 1808 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_13
timestamp 1524952243
transform -1 0 1920 0 1 1170
box -8 -3 64 105
use NAND2X1  NAND2X1_21
timestamp 1524952243
transform -1 0 1944 0 1 1170
box -8 -3 32 105
use top_module_VIA0  top_module_VIA0_15
timestamp 1524952243
transform 1 0 1970 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_885
timestamp 1524952243
transform 1 0 68 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1524952243
transform 1 0 132 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1524952243
transform 1 0 172 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_926
timestamp 1524952243
transform 1 0 156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1524952243
transform 1 0 172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1524952243
transform 1 0 76 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_951
timestamp 1524952243
transform 1 0 124 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_987
timestamp 1524952243
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_876
timestamp 1524952243
transform 1 0 244 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1524952243
transform 1 0 204 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1524952243
transform 1 0 228 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1524952243
transform 1 0 252 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1524952243
transform 1 0 196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1524952243
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1524952243
transform 1 0 188 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1046
timestamp 1524952243
transform 1 0 172 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_941
timestamp 1524952243
transform 1 0 212 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_930
timestamp 1524952243
transform 1 0 300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1524952243
transform 1 0 316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1524952243
transform 1 0 212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1524952243
transform 1 0 220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1524952243
transform 1 0 276 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_913
timestamp 1524952243
transform 1 0 324 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1524952243
transform 1 0 340 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1524952243
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1524952243
transform 1 0 356 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_953
timestamp 1524952243
transform 1 0 324 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1524952243
transform 1 0 340 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_972
timestamp 1524952243
transform 1 0 276 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1524952243
transform 1 0 316 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1524952243
transform 1 0 356 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_924
timestamp 1524952243
transform 1 0 388 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1524952243
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_942
timestamp 1524952243
transform 1 0 388 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1524952243
transform 1 0 372 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1524952243
transform 1 0 324 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_995
timestamp 1524952243
transform 1 0 220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1524952243
transform 1 0 300 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1524952243
transform 1 0 348 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_1048
timestamp 1524952243
transform 1 0 356 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_996
timestamp 1524952243
transform 1 0 356 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1524952243
transform 1 0 412 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_935
timestamp 1524952243
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_943
timestamp 1524952243
transform 1 0 428 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_936
timestamp 1524952243
transform 1 0 436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1524952243
transform 1 0 404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1524952243
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1524952243
transform 1 0 428 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_975
timestamp 1524952243
transform 1 0 412 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_1049
timestamp 1524952243
transform 1 0 428 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_997
timestamp 1524952243
transform 1 0 428 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1524952243
transform 1 0 484 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1524952243
transform 1 0 468 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_937
timestamp 1524952243
transform 1 0 476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1524952243
transform 1 0 484 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_877
timestamp 1524952243
transform 1 0 500 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1524952243
transform 1 0 508 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_996
timestamp 1524952243
transform 1 0 460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1524952243
transform 1 0 484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1524952243
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1524952243
transform 1 0 460 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_976
timestamp 1524952243
transform 1 0 484 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1524952243
transform 1 0 460 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1524952243
transform 1 0 508 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1051
timestamp 1524952243
transform 1 0 500 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1524952243
transform 1 0 524 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_939
timestamp 1524952243
transform 1 0 532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1524952243
transform 1 0 524 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_956
timestamp 1524952243
transform 1 0 532 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1052
timestamp 1524952243
transform 1 0 532 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1524952243
transform 1 0 524 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1524952243
transform 1 0 516 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1524952243
transform 1 0 556 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1524952243
transform 1 0 612 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1524952243
transform 1 0 644 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1524952243
transform 1 0 676 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1524952243
transform 1 0 604 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_940
timestamp 1524952243
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1524952243
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1524952243
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1524952243
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1524952243
transform 1 0 604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1524952243
transform 1 0 644 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_1017
timestamp 1524952243
transform 1 0 548 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1524952243
transform 1 0 652 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1524952243
transform 1 0 588 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1524952243
transform 1 0 644 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1524952243
transform 1 0 684 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1524952243
transform 1 0 700 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_943
timestamp 1524952243
transform 1 0 684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1524952243
transform 1 0 700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1524952243
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1524952243
transform 1 0 676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1524952243
transform 1 0 692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_958
timestamp 1524952243
transform 1 0 700 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1524952243
transform 1 0 740 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_946
timestamp 1524952243
transform 1 0 724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1524952243
transform 1 0 748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1524952243
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1524952243
transform 1 0 732 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_977
timestamp 1524952243
transform 1 0 708 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1524952243
transform 1 0 700 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1524952243
transform 1 0 740 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1524952243
transform 1 0 772 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1524952243
transform 1 0 788 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1524952243
transform 1 0 780 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_945
timestamp 1524952243
transform 1 0 788 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_1007
timestamp 1524952243
transform 1 0 772 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1524952243
transform 1 0 756 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1524952243
transform 1 0 812 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1524952243
transform 1 0 804 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_1008
timestamp 1524952243
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1524952243
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1524952243
transform 1 0 804 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1524952243
transform 1 0 796 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1524952243
transform 1 0 972 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1524952243
transform 1 0 868 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1524952243
transform 1 0 908 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_949
timestamp 1524952243
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1524952243
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_947
timestamp 1524952243
transform 1 0 852 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_951
timestamp 1524952243
transform 1 0 868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1524952243
transform 1 0 884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1524952243
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_959
timestamp 1524952243
transform 1 0 836 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1524952243
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1524952243
transform 1 0 836 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1524952243
transform 1 0 868 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1524952243
transform 1 0 884 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1524952243
transform 1 0 908 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1524952243
transform 1 0 964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1524952243
transform 1 0 868 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1524952243
transform 1 0 1108 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1524952243
transform 1 0 1148 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1524952243
transform 1 0 1164 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1524952243
transform 1 0 1132 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1524952243
transform 1 0 1196 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1524952243
transform 1 0 1228 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1524952243
transform 1 0 1268 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1524952243
transform 1 0 1292 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1524952243
transform 1 0 1172 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1524952243
transform 1 0 1188 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1524952243
transform 1 0 1212 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_954
timestamp 1524952243
transform 1 0 996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1524952243
transform 1 0 1012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1524952243
transform 1 0 1100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1524952243
transform 1 0 1116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1524952243
transform 1 0 1132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1524952243
transform 1 0 1140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1524952243
transform 1 0 1156 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_962
timestamp 1524952243
transform 1 0 980 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1013
timestamp 1524952243
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1524952243
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1524952243
transform 1 0 972 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_1000
timestamp 1524952243
transform 1 0 844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1524952243
transform 1 0 868 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1524952243
transform 1 0 900 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1524952243
transform 1 0 860 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1524952243
transform 1 0 836 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1524952243
transform 1 0 924 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1524952243
transform 1 0 956 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1524952243
transform 1 0 964 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1524952243
transform 1 0 1060 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1524952243
transform 1 0 1100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1524952243
transform 1 0 1108 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1524952243
transform 1 0 1116 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1524952243
transform 1 0 1124 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_948
timestamp 1524952243
transform 1 0 1164 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1524952243
transform 1 0 1324 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1524952243
transform 1 0 1316 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1524952243
transform 1 0 1364 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1524952243
transform 1 0 1508 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1524952243
transform 1 0 1468 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1524952243
transform 1 0 1500 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1524952243
transform 1 0 1348 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1524952243
transform 1 0 1380 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1524952243
transform 1 0 1452 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_961
timestamp 1524952243
transform 1 0 1172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1524952243
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1524952243
transform 1 0 1196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1524952243
transform 1 0 1212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1524952243
transform 1 0 1228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1524952243
transform 1 0 1316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1524952243
transform 1 0 1340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1524952243
transform 1 0 1148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1524952243
transform 1 0 1164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1524952243
transform 1 0 1180 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_965
timestamp 1524952243
transform 1 0 1188 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1524952243
transform 1 0 1204 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_980
timestamp 1524952243
transform 1 0 1132 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1524952243
transform 1 0 1148 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1524952243
transform 1 0 1180 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1524952243
transform 1 0 1196 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1524952243
transform 1 0 1108 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1524952243
transform 1 0 1100 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1524952243
transform 1 0 1180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1524952243
transform 1 0 1196 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_968
timestamp 1524952243
transform 1 0 1364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1524952243
transform 1 0 1452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1524952243
transform 1 0 1252 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1524952243
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1524952243
transform 1 0 1316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1524952243
transform 1 0 1332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1524952243
transform 1 0 1348 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_984
timestamp 1524952243
transform 1 0 1252 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1524952243
transform 1 0 1308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1524952243
transform 1 0 1244 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1524952243
transform 1 0 1380 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1524952243
transform 1 0 1388 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_1007
timestamp 1524952243
transform 1 0 1412 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1524952243
transform 1 0 1508 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1524952243
transform 1 0 1556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1524952243
transform 1 0 1596 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1524952243
transform 1 0 1628 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1524952243
transform 1 0 1540 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_970
timestamp 1524952243
transform 1 0 1508 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_949
timestamp 1524952243
transform 1 0 1516 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1524952243
transform 1 0 1532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1524952243
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1524952243
transform 1 0 1508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1524952243
transform 1 0 1524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1524952243
transform 1 0 1540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1524952243
transform 1 0 1548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_986
timestamp 1524952243
transform 1 0 1532 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1524952243
transform 1 0 1476 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1524952243
transform 1 0 1508 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1524952243
transform 1 0 1444 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1524952243
transform 1 0 1388 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1524952243
transform 1 0 1548 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1524952243
transform 1 0 1532 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1524952243
transform 1 0 1604 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1524952243
transform 1 0 1604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1524952243
transform 1 0 1612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1524952243
transform 1 0 1628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1524952243
transform 1 0 1636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1524952243
transform 1 0 1604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1524952243
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_967
timestamp 1524952243
transform 1 0 1628 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1524952243
transform 1 0 1700 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1524952243
transform 1 0 1716 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1524952243
transform 1 0 1732 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1524952243
transform 1 0 1692 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_976
timestamp 1524952243
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1524952243
transform 1 0 1700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1524952243
transform 1 0 1644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1524952243
transform 1 0 1676 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_968
timestamp 1524952243
transform 1 0 1692 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1524952243
transform 1 0 1732 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1524952243
transform 1 0 1780 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1524952243
transform 1 0 1764 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1524952243
transform 1 0 1812 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1524952243
transform 1 0 1844 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_978
timestamp 1524952243
transform 1 0 1764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1524952243
transform 1 0 1780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1524952243
transform 1 0 1796 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1524952243
transform 1 0 1748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1524952243
transform 1 0 1756 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_987
timestamp 1524952243
transform 1 0 1612 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1524952243
transform 1 0 1644 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1524952243
transform 1 0 1676 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1524952243
transform 1 0 1604 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1524952243
transform 1 0 1556 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1524952243
transform 1 0 1636 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1524952243
transform 1 0 1764 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1039
timestamp 1524952243
transform 1 0 1772 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1524952243
transform 1 0 1788 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_990
timestamp 1524952243
transform 1 0 1748 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1524952243
transform 1 0 1788 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1524952243
transform 1 0 1780 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1524952243
transform 1 0 1916 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1524952243
transform 1 0 1924 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1524952243
transform 1 0 1876 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1524952243
transform 1 0 1892 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1524952243
transform 1 0 1844 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1524952243
transform 1 0 1852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1524952243
transform 1 0 1860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1524952243
transform 1 0 1876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1524952243
transform 1 0 1892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1524952243
transform 1 0 1940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1524952243
transform 1 0 1844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1524952243
transform 1 0 1852 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_971
timestamp 1524952243
transform 1 0 1860 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1524952243
transform 1 0 1868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1524952243
transform 1 0 1884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1524952243
transform 1 0 1908 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_992
timestamp 1524952243
transform 1 0 1844 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1524952243
transform 1 0 1884 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1524952243
transform 1 0 1908 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1524952243
transform 1 0 1876 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1524952243
transform 1 0 1924 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1524952243
transform 1 0 1900 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1524952243
transform 1 0 1940 0 1 1085
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_16
timestamp 1524952243
transform 1 0 24 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_1035
timestamp 1524952243
transform 1 0 76 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1524952243
transform 1 0 172 0 1 1075
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_48
timestamp 1524952243
transform -1 0 168 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_40
timestamp 1524952243
transform -1 0 200 0 -1 1170
box -8 -3 34 105
use INVX2  INVX2_71
timestamp 1524952243
transform 1 0 200 0 -1 1170
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_53
timestamp 1524952243
transform -1 0 312 0 -1 1170
box -8 -3 104 105
use FILL  FILL_13
timestamp 1524952243
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_41
timestamp 1524952243
transform -1 0 352 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1524952243
transform -1 0 384 0 -1 1170
box -8 -3 34 105
use NOR2X1  NOR2X1_25
timestamp 1524952243
transform 1 0 384 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1524952243
transform 1 0 408 0 -1 1170
box -8 -3 32 105
use BUFX2  BUFX2_7
timestamp 1524952243
transform -1 0 456 0 -1 1170
box -5 -3 28 105
use NAND2X1  NAND2X1_23
timestamp 1524952243
transform -1 0 480 0 -1 1170
box -8 -3 32 105
use M3_M2  M3_M2_1037
timestamp 1524952243
transform 1 0 492 0 1 1075
box -3 -3 3 3
use NAND2X1  NAND2X1_24
timestamp 1524952243
transform 1 0 480 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1524952243
transform -1 0 528 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1524952243
transform -1 0 552 0 -1 1170
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_54
timestamp 1524952243
transform 1 0 552 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_72
timestamp 1524952243
transform 1 0 648 0 -1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_3
timestamp 1524952243
transform 1 0 664 0 -1 1170
box -8 -3 46 105
use INVX2  INVX2_73
timestamp 1524952243
transform 1 0 704 0 -1 1170
box -9 -3 26 105
use M3_M2  M3_M2_1038
timestamp 1524952243
transform 1 0 740 0 1 1075
box -3 -3 3 3
use OAI21X1  OAI21X1_43
timestamp 1524952243
transform 1 0 720 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1524952243
transform -1 0 784 0 -1 1170
box -8 -3 34 105
use M3_M2  M3_M2_1039
timestamp 1524952243
transform 1 0 812 0 1 1075
box -3 -3 3 3
use NOR2X1  NOR2X1_26
timestamp 1524952243
transform 1 0 784 0 -1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_45
timestamp 1524952243
transform 1 0 808 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1524952243
transform 1 0 840 0 -1 1170
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_55
timestamp 1524952243
transform 1 0 872 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_47
timestamp 1524952243
transform -1 0 1000 0 -1 1170
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_56
timestamp 1524952243
transform 1 0 1000 0 -1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_4
timestamp 1524952243
transform 1 0 1096 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1524952243
transform 1 0 1136 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1524952243
transform 1 0 1176 0 -1 1170
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_57
timestamp 1524952243
transform 1 0 1216 0 -1 1170
box -8 -3 104 105
use AOI22X1  AOI22X1_22
timestamp 1524952243
transform 1 0 1312 0 -1 1170
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_58
timestamp 1524952243
transform 1 0 1352 0 -1 1170
box -8 -3 104 105
use M3_M2  M3_M2_1040
timestamp 1524952243
transform 1 0 1508 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1524952243
transform 1 0 1524 0 1 1075
box -3 -3 3 3
use XOR2X1  XOR2X1_14
timestamp 1524952243
transform 1 0 1448 0 -1 1170
box -8 -3 64 105
use AOI22X1  AOI22X1_23
timestamp 1524952243
transform -1 0 1544 0 -1 1170
box -8 -3 46 105
use XNOR2X1  XNOR2X1_8
timestamp 1524952243
transform -1 0 1600 0 -1 1170
box -8 -3 64 105
use AOI22X1  AOI22X1_24
timestamp 1524952243
transform 1 0 1600 0 -1 1170
box -8 -3 46 105
use XNOR2X1  XNOR2X1_9
timestamp 1524952243
transform 1 0 1640 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_10
timestamp 1524952243
transform 1 0 1696 0 -1 1170
box -8 -3 64 105
use M3_M2  M3_M2_1042
timestamp 1524952243
transform 1 0 1788 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_25
timestamp 1524952243
transform -1 0 1792 0 -1 1170
box -8 -3 46 105
use XNOR2X1  XNOR2X1_11
timestamp 1524952243
transform 1 0 1792 0 -1 1170
box -8 -3 64 105
use AOI22X1  AOI22X1_26
timestamp 1524952243
transform 1 0 1848 0 -1 1170
box -8 -3 46 105
use XOR2X1  XOR2X1_15
timestamp 1524952243
transform -1 0 1944 0 -1 1170
box -8 -3 64 105
use top_module_VIA0  top_module_VIA0_17
timestamp 1524952243
transform 1 0 1994 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_1082
timestamp 1524952243
transform 1 0 76 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1073
timestamp 1524952243
transform 1 0 68 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1118
timestamp 1524952243
transform 1 0 116 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1524952243
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1119
timestamp 1524952243
transform 1 0 156 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1058
timestamp 1524952243
transform 1 0 188 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1524952243
transform 1 0 156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1524952243
transform 1 0 172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1524952243
transform 1 0 188 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1162
timestamp 1524952243
transform 1 0 132 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1524952243
transform 1 0 76 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1524952243
transform 1 0 204 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1524952243
transform 1 0 220 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1059
timestamp 1524952243
transform 1 0 228 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1524952243
transform 1 0 212 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1163
timestamp 1524952243
transform 1 0 188 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_1076
timestamp 1524952243
transform 1 0 236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1524952243
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1164
timestamp 1524952243
transform 1 0 228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1524952243
transform 1 0 212 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1524952243
transform 1 0 276 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1060
timestamp 1524952243
transform 1 0 268 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_1120
timestamp 1524952243
transform 1 0 260 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1077
timestamp 1524952243
transform 1 0 268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1524952243
transform 1 0 276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1524952243
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1524952243
transform 1 0 300 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1524952243
transform 1 0 292 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1524952243
transform 1 0 300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1524952243
transform 1 0 284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1524952243
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1141
timestamp 1524952243
transform 1 0 300 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1142
timestamp 1524952243
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1165
timestamp 1524952243
transform 1 0 284 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_1202
timestamp 1524952243
transform 1 0 300 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_1142
timestamp 1524952243
transform 1 0 316 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1143
timestamp 1524952243
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1056
timestamp 1524952243
transform 1 0 340 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1524952243
transform 1 0 388 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1524952243
transform 1 0 420 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1524952243
transform 1 0 348 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1524952243
transform 1 0 372 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1524952243
transform 1 0 396 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1524952243
transform 1 0 468 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1524952243
transform 1 0 356 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1080
timestamp 1524952243
transform 1 0 332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1524952243
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1524952243
transform 1 0 332 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1524952243
transform 1 0 436 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1082
timestamp 1524952243
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1524952243
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1524952243
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1524952243
transform 1 0 356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1524952243
transform 1 0 364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1524952243
transform 1 0 388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1524952243
transform 1 0 404 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1524952243
transform 1 0 316 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1524952243
transform 1 0 324 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1524952243
transform 1 0 316 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1524952243
transform 1 0 340 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1524952243
transform 1 0 428 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1524952243
transform 1 0 596 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1524952243
transform 1 0 548 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1524952243
transform 1 0 596 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1524952243
transform 1 0 644 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1524952243
transform 1 0 708 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1524952243
transform 1 0 724 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1524952243
transform 1 0 700 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1524952243
transform 1 0 644 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1085
timestamp 1524952243
transform 1 0 500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1524952243
transform 1 0 556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1524952243
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1524952243
transform 1 0 612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1524952243
transform 1 0 628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1524952243
transform 1 0 644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1524952243
transform 1 0 492 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1524952243
transform 1 0 372 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1524952243
transform 1 0 388 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1524952243
transform 1 0 500 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1149
timestamp 1524952243
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1169
timestamp 1524952243
transform 1 0 492 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1524952243
transform 1 0 380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1524952243
transform 1 0 396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1524952243
transform 1 0 452 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1524952243
transform 1 0 596 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1150
timestamp 1524952243
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1524952243
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1524952243
transform 1 0 628 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1524952243
transform 1 0 676 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1091
timestamp 1524952243
transform 1 0 700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1524952243
transform 1 0 636 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1170
timestamp 1524952243
transform 1 0 556 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1524952243
transform 1 0 684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1524952243
transform 1 0 700 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1524952243
transform 1 0 756 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1524952243
transform 1 0 772 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_1061
timestamp 1524952243
transform 1 0 764 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1524952243
transform 1 0 772 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1092
timestamp 1524952243
transform 1 0 748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1524952243
transform 1 0 764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1524952243
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1524952243
transform 1 0 740 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1171
timestamp 1524952243
transform 1 0 620 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1524952243
transform 1 0 644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1524952243
transform 1 0 676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1524952243
transform 1 0 700 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1524952243
transform 1 0 756 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1155
timestamp 1524952243
transform 1 0 764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1524952243
transform 1 0 772 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1524952243
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1524952243
transform 1 0 788 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1204
timestamp 1524952243
transform 1 0 788 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1524952243
transform 1 0 836 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1524952243
transform 1 0 828 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1524952243
transform 1 0 836 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1062
timestamp 1524952243
transform 1 0 844 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1524952243
transform 1 0 812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1524952243
transform 1 0 828 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1191
timestamp 1524952243
transform 1 0 788 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1524952243
transform 1 0 804 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1524952243
transform 1 0 908 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1524952243
transform 1 0 876 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1524952243
transform 1 0 892 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1524952243
transform 1 0 924 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1524952243
transform 1 0 860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1524952243
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1524952243
transform 1 0 844 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1524952243
transform 1 0 852 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1152
timestamp 1524952243
transform 1 0 860 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1098
timestamp 1524952243
transform 1 0 884 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1524952243
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1524952243
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1524952243
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1524952243
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1524952243
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1524952243
transform 1 0 916 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1100
timestamp 1524952243
transform 1 0 948 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1101
timestamp 1524952243
transform 1 0 940 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1193
timestamp 1524952243
transform 1 0 916 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1524952243
transform 1 0 956 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1524952243
transform 1 0 980 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1524952243
transform 1 0 1004 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1524952243
transform 1 0 1028 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1524952243
transform 1 0 1044 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_1057
timestamp 1524952243
transform 1 0 1044 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_1091
timestamp 1524952243
transform 1 0 1060 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1524952243
transform 1 0 1100 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1524952243
transform 1 0 980 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1524952243
transform 1 0 988 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1524952243
transform 1 0 1004 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1524952243
transform 1 0 1028 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1524952243
transform 1 0 964 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1124
timestamp 1524952243
transform 1 0 988 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1524952243
transform 1 0 996 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1524952243
transform 1 0 948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1524952243
transform 1 0 956 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1153
timestamp 1524952243
transform 1 0 972 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1166
timestamp 1524952243
transform 1 0 980 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1154
timestamp 1524952243
transform 1 0 988 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1524952243
transform 1 0 1044 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1068
timestamp 1524952243
transform 1 0 1052 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1524952243
transform 1 0 1076 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1524952243
transform 1 0 1028 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1104
timestamp 1524952243
transform 1 0 1036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1524952243
transform 1 0 1012 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1194
timestamp 1524952243
transform 1 0 956 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1524952243
transform 1 0 988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1524952243
transform 1 0 1012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1524952243
transform 1 0 1052 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1105
timestamp 1524952243
transform 1 0 1060 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1048
timestamp 1524952243
transform 1 0 1156 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1524952243
transform 1 0 1180 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1524952243
transform 1 0 1148 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1524952243
transform 1 0 1156 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1524952243
transform 1 0 1140 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1524952243
transform 1 0 1164 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1069
timestamp 1524952243
transform 1 0 1172 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1524952243
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1127
timestamp 1524952243
transform 1 0 1108 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1524952243
transform 1 0 1124 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1107
timestamp 1524952243
transform 1 0 1132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1524952243
transform 1 0 1140 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1129
timestamp 1524952243
transform 1 0 1148 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1524952243
transform 1 0 1212 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1524952243
transform 1 0 1244 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_1070
timestamp 1524952243
transform 1 0 1204 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_1105
timestamp 1524952243
transform 1 0 1220 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1524952243
transform 1 0 1300 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1524952243
transform 1 0 1260 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_1071
timestamp 1524952243
transform 1 0 1236 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1524952243
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1524952243
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1524952243
transform 1 0 1188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1524952243
transform 1 0 1068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1524952243
transform 1 0 1076 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1197
timestamp 1524952243
transform 1 0 1052 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1524952243
transform 1 0 1124 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1524952243
transform 1 0 1132 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1171
timestamp 1524952243
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1524952243
transform 1 0 1148 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1198
timestamp 1524952243
transform 1 0 1124 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1524952243
transform 1 0 1204 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1524952243
transform 1 0 1252 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1072
timestamp 1524952243
transform 1 0 1260 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1524952243
transform 1 0 1212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1524952243
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1524952243
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1524952243
transform 1 0 1188 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1524952243
transform 1 0 1236 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1175
timestamp 1524952243
transform 1 0 1204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1524952243
transform 1 0 1212 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1157
timestamp 1524952243
transform 1 0 1228 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1177
timestamp 1524952243
transform 1 0 1236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1524952243
transform 1 0 1244 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1199
timestamp 1524952243
transform 1 0 1204 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1524952243
transform 1 0 1252 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1524952243
transform 1 0 1284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1524952243
transform 1 0 1300 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1524952243
transform 1 0 1380 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1524952243
transform 1 0 1388 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1113
timestamp 1524952243
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1524952243
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1524952243
transform 1 0 1380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1524952243
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1524952243
transform 1 0 1260 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_1180
timestamp 1524952243
transform 1 0 1316 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1524952243
transform 1 0 1316 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1524952243
transform 1 0 1268 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1524952243
transform 1 0 1284 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1524952243
transform 1 0 1300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1524952243
transform 1 0 1396 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1524952243
transform 1 0 1444 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1524952243
transform 1 0 1508 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1524952243
transform 1 0 1524 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1524952243
transform 1 0 1540 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1524952243
transform 1 0 1500 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1116
timestamp 1524952243
transform 1 0 1428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1524952243
transform 1 0 1444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1524952243
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1524952243
transform 1 0 1372 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1159
timestamp 1524952243
transform 1 0 1380 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1524952243
transform 1 0 1388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1524952243
transform 1 0 1396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1203
timestamp 1524952243
transform 1 0 1364 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1524952243
transform 1 0 1380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1524952243
transform 1 0 1484 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1524952243
transform 1 0 1588 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1524952243
transform 1 0 1612 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1524952243
transform 1 0 1556 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1524952243
transform 1 0 1580 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1119
timestamp 1524952243
transform 1 0 1500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1524952243
transform 1 0 1508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1524952243
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1135
timestamp 1524952243
transform 1 0 1524 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1121
timestamp 1524952243
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1524952243
transform 1 0 1572 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1524952243
transform 1 0 1580 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1137
timestamp 1524952243
transform 1 0 1588 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1524952243
transform 1 0 1636 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1123
timestamp 1524952243
transform 1 0 1596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1524952243
transform 1 0 1612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1524952243
transform 1 0 1628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1524952243
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1160
timestamp 1524952243
transform 1 0 1500 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1185
timestamp 1524952243
transform 1 0 1508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1524952243
transform 1 0 1524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1524952243
transform 1 0 1580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1524952243
transform 1 0 1588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1524952243
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1524952243
transform 1 0 1620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1524952243
transform 1 0 1636 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1177
timestamp 1524952243
transform 1 0 1636 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1524952243
transform 1 0 1612 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1524952243
transform 1 0 1700 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1524952243
transform 1 0 1684 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1524952243
transform 1 0 1708 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1524952243
transform 1 0 1684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1524952243
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1524952243
transform 1 0 1684 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1178
timestamp 1524952243
transform 1 0 1684 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1524952243
transform 1 0 1676 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1524952243
transform 1 0 1772 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1524952243
transform 1 0 1796 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1524952243
transform 1 0 1780 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1524952243
transform 1 0 1756 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1129
timestamp 1524952243
transform 1 0 1764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1524952243
transform 1 0 1780 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1524952243
transform 1 0 1748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1524952243
transform 1 0 1756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1524952243
transform 1 0 1788 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1179
timestamp 1524952243
transform 1 0 1740 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1524952243
transform 1 0 1756 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1524952243
transform 1 0 1772 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1524952243
transform 1 0 1836 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_1131
timestamp 1524952243
transform 1 0 1844 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_1140
timestamp 1524952243
transform 1 0 1860 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1524952243
transform 1 0 1908 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1524952243
transform 1 0 1932 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1524952243
transform 1 0 1916 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1524952243
transform 1 0 1948 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1524952243
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1524952243
transform 1 0 1916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1524952243
transform 1 0 1932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1524952243
transform 1 0 1836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1524952243
transform 1 0 1844 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1161
timestamp 1524952243
transform 1 0 1892 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_1198
timestamp 1524952243
transform 1 0 1900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1524952243
transform 1 0 1908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1524952243
transform 1 0 1924 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1182
timestamp 1524952243
transform 1 0 1844 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_1201
timestamp 1524952243
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_1183
timestamp 1524952243
transform 1 0 1932 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1524952243
transform 1 0 1892 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1524952243
transform 1 0 1916 0 1 985
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_18
timestamp 1524952243
transform 1 0 48 0 1 970
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_59
timestamp 1524952243
transform -1 0 168 0 1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_27
timestamp 1524952243
transform 1 0 168 0 1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_48
timestamp 1524952243
transform -1 0 224 0 1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_28
timestamp 1524952243
transform -1 0 248 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_1209
timestamp 1524952243
transform 1 0 268 0 1 975
box -3 -3 3 3
use NAND2X1  NAND2X1_29
timestamp 1524952243
transform 1 0 248 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1524952243
transform -1 0 296 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1524952243
transform -1 0 320 0 1 970
box -8 -3 32 105
use INVX2  INVX2_74
timestamp 1524952243
transform 1 0 320 0 1 970
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1524952243
transform -1 0 352 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_27
timestamp 1524952243
transform -1 0 392 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_1210
timestamp 1524952243
transform 1 0 420 0 1 975
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_60
timestamp 1524952243
transform 1 0 392 0 1 970
box -8 -3 104 105
use INVX2  INVX2_76
timestamp 1524952243
transform 1 0 488 0 1 970
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_61
timestamp 1524952243
transform 1 0 504 0 1 970
box -8 -3 104 105
use OAI22X1  OAI22X1_7
timestamp 1524952243
transform 1 0 600 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_1211
timestamp 1524952243
transform 1 0 684 0 1 975
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_62
timestamp 1524952243
transform -1 0 736 0 1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_49
timestamp 1524952243
transform 1 0 736 0 1 970
box -8 -3 34 105
use NOR2X1  NOR2X1_29
timestamp 1524952243
transform -1 0 792 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1524952243
transform 1 0 792 0 1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_50
timestamp 1524952243
transform 1 0 816 0 1 970
box -8 -3 34 105
use INVX2  INVX2_77
timestamp 1524952243
transform 1 0 848 0 1 970
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1524952243
transform -1 0 880 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_28
timestamp 1524952243
transform 1 0 880 0 1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_51
timestamp 1524952243
transform -1 0 952 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1524952243
transform 1 0 952 0 1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_30
timestamp 1524952243
transform -1 0 1008 0 1 970
box -8 -3 32 105
use INVX2  INVX2_79
timestamp 1524952243
transform 1 0 1008 0 1 970
box -9 -3 26 105
use NAND3X1  NAND3X1_17
timestamp 1524952243
transform 1 0 1024 0 1 970
box -8 -3 40 105
use INVX2  INVX2_80
timestamp 1524952243
transform -1 0 1072 0 1 970
box -9 -3 26 105
use XOR2X1  XOR2X1_16
timestamp 1524952243
transform 1 0 1072 0 1 970
box -8 -3 64 105
use INVX2  INVX2_81
timestamp 1524952243
transform -1 0 1144 0 1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_53
timestamp 1524952243
transform 1 0 1144 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1524952243
transform 1 0 1176 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1524952243
transform 1 0 1208 0 1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_31
timestamp 1524952243
transform 1 0 1240 0 1 970
box -8 -3 32 105
use XOR2X1  XOR2X1_17
timestamp 1524952243
transform 1 0 1264 0 1 970
box -8 -3 64 105
use M3_M2  M3_M2_1212
timestamp 1524952243
transform 1 0 1372 0 1 975
box -3 -3 3 3
use XNOR2X1  XNOR2X1_12
timestamp 1524952243
transform 1 0 1320 0 1 970
box -8 -3 64 105
use INVX2  INVX2_82
timestamp 1524952243
transform -1 0 1392 0 1 970
box -9 -3 26 105
use XOR2X1  XOR2X1_18
timestamp 1524952243
transform 1 0 1392 0 1 970
box -8 -3 64 105
use M3_M2  M3_M2_1213
timestamp 1524952243
transform 1 0 1508 0 1 975
box -3 -3 3 3
use XNOR2X1  XNOR2X1_13
timestamp 1524952243
transform -1 0 1504 0 1 970
box -8 -3 64 105
use INVX2  INVX2_83
timestamp 1524952243
transform 1 0 1504 0 1 970
box -9 -3 26 105
use XOR2X1  XOR2X1_19
timestamp 1524952243
transform 1 0 1520 0 1 970
box -8 -3 64 105
use AOI22X1  AOI22X1_29
timestamp 1524952243
transform -1 0 1616 0 1 970
box -8 -3 46 105
use INVX2  INVX2_84
timestamp 1524952243
transform 1 0 1616 0 1 970
box -9 -3 26 105
use XNOR2X1  XNOR2X1_14
timestamp 1524952243
transform -1 0 1688 0 1 970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_15
timestamp 1524952243
transform -1 0 1744 0 1 970
box -8 -3 64 105
use AOI22X1  AOI22X1_30
timestamp 1524952243
transform 1 0 1744 0 1 970
box -8 -3 46 105
use XOR2X1  XOR2X1_20
timestamp 1524952243
transform 1 0 1784 0 1 970
box -8 -3 64 105
use M3_M2  M3_M2_1214
timestamp 1524952243
transform 1 0 1860 0 1 975
box -3 -3 3 3
use XNOR2X1  XNOR2X1_16
timestamp 1524952243
transform 1 0 1840 0 1 970
box -8 -3 64 105
use M3_M2  M3_M2_1215
timestamp 1524952243
transform 1 0 1908 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_31
timestamp 1524952243
transform -1 0 1936 0 1 970
box -8 -3 46 105
use FILL  FILL_14
timestamp 1524952243
transform 1 0 1936 0 1 970
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_19
timestamp 1524952243
transform 1 0 1970 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_1216
timestamp 1524952243
transform 1 0 140 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1524952243
transform 1 0 76 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1524952243
transform 1 0 156 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1524952243
transform 1 0 124 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1524952243
transform 1 0 172 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1524952243
transform 1 0 196 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1524952243
transform 1 0 132 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1210
timestamp 1524952243
transform 1 0 156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1524952243
transform 1 0 172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1524952243
transform 1 0 196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1524952243
transform 1 0 76 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1524952243
transform 1 0 132 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1327
timestamp 1524952243
transform 1 0 76 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_1266
timestamp 1524952243
transform 1 0 188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1524952243
transform 1 0 196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1524952243
transform 1 0 172 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1217
timestamp 1524952243
transform 1 0 228 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1524952243
transform 1 0 236 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1524952243
transform 1 0 276 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1524952243
transform 1 0 228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1524952243
transform 1 0 236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1524952243
transform 1 0 220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1524952243
transform 1 0 204 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1342
timestamp 1524952243
transform 1 0 172 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1524952243
transform 1 0 196 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1524952243
transform 1 0 220 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1524952243
transform 1 0 140 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1524952243
transform 1 0 188 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1524952243
transform 1 0 244 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1215
timestamp 1524952243
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1524952243
transform 1 0 276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1524952243
transform 1 0 244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1378
timestamp 1524952243
transform 1 0 236 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1524952243
transform 1 0 252 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1524952243
transform 1 0 284 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1524952243
transform 1 0 316 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1524952243
transform 1 0 316 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1524952243
transform 1 0 316 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1270
timestamp 1524952243
transform 1 0 268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1524952243
transform 1 0 284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1303
timestamp 1524952243
transform 1 0 292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1272
timestamp 1524952243
transform 1 0 300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1524952243
transform 1 0 252 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1328
timestamp 1524952243
transform 1 0 276 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_1337
timestamp 1524952243
transform 1 0 284 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1345
timestamp 1524952243
transform 1 0 300 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1524952243
transform 1 0 268 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1524952243
transform 1 0 284 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1524952243
transform 1 0 316 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1524952243
transform 1 0 332 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1217
timestamp 1524952243
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1524952243
transform 1 0 332 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1236
timestamp 1524952243
transform 1 0 404 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1524952243
transform 1 0 420 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1524952243
transform 1 0 444 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1524952243
transform 1 0 364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1524952243
transform 1 0 380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1524952243
transform 1 0 388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1524952243
transform 1 0 356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1524952243
transform 1 0 372 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1304
timestamp 1524952243
transform 1 0 380 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1524952243
transform 1 0 404 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1221
timestamp 1524952243
transform 1 0 420 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1288
timestamp 1524952243
transform 1 0 468 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1276
timestamp 1524952243
transform 1 0 388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1524952243
transform 1 0 404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1524952243
transform 1 0 444 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1329
timestamp 1524952243
transform 1 0 364 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1524952243
transform 1 0 348 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1524952243
transform 1 0 372 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1524952243
transform 1 0 492 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1524952243
transform 1 0 532 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1524952243
transform 1 0 572 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1524952243
transform 1 0 516 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1524952243
transform 1 0 636 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1222
timestamp 1524952243
transform 1 0 532 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1524952243
transform 1 0 612 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1524952243
transform 1 0 724 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1524952243
transform 1 0 668 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1223
timestamp 1524952243
transform 1 0 620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1524952243
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1524952243
transform 1 0 652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1524952243
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1524952243
transform 1 0 500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1524952243
transform 1 0 516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1524952243
transform 1 0 572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1524952243
transform 1 0 612 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1330
timestamp 1524952243
transform 1 0 404 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1524952243
transform 1 0 444 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1524952243
transform 1 0 420 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1524952243
transform 1 0 484 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1524952243
transform 1 0 436 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1524952243
transform 1 0 620 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1283
timestamp 1524952243
transform 1 0 628 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1307
timestamp 1524952243
transform 1 0 636 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1284
timestamp 1524952243
transform 1 0 644 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1291
timestamp 1524952243
transform 1 0 692 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1524952243
transform 1 0 732 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1524952243
transform 1 0 796 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1524952243
transform 1 0 820 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1524952243
transform 1 0 772 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1524952243
transform 1 0 780 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1524952243
transform 1 0 820 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1524952243
transform 1 0 868 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1227
timestamp 1524952243
transform 1 0 756 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1293
timestamp 1524952243
transform 1 0 764 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1228
timestamp 1524952243
transform 1 0 780 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1294
timestamp 1524952243
transform 1 0 812 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1285
timestamp 1524952243
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1524952243
transform 1 0 756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1524952243
transform 1 0 764 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1308
timestamp 1524952243
transform 1 0 780 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1288
timestamp 1524952243
transform 1 0 820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1524952243
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1524952243
transform 1 0 868 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1332
timestamp 1524952243
transform 1 0 684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1524952243
transform 1 0 748 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1524952243
transform 1 0 628 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1524952243
transform 1 0 652 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1524952243
transform 1 0 876 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_1229
timestamp 1524952243
transform 1 0 876 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1524952243
transform 1 0 884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1524952243
transform 1 0 876 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1223
timestamp 1524952243
transform 1 0 956 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1524952243
transform 1 0 948 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1206
timestamp 1524952243
transform 1 0 900 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_1267
timestamp 1524952243
transform 1 0 908 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1524952243
transform 1 0 932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1524952243
transform 1 0 900 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1231
timestamp 1524952243
transform 1 0 908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1524952243
transform 1 0 932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1524952243
transform 1 0 892 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1296
timestamp 1524952243
transform 1 0 940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1524952243
transform 1 0 1004 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1524952243
transform 1 0 1020 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1524952243
transform 1 0 980 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1524952243
transform 1 0 964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1524952243
transform 1 0 924 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1524952243
transform 1 0 940 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1309
timestamp 1524952243
transform 1 0 956 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1295
timestamp 1524952243
transform 1 0 964 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1334
timestamp 1524952243
transform 1 0 940 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_1338
timestamp 1524952243
transform 1 0 956 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1351
timestamp 1524952243
transform 1 0 956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1524952243
transform 1 0 948 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1524952243
transform 1 0 980 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1524952243
transform 1 0 1068 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1524952243
transform 1 0 1052 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1234
timestamp 1524952243
transform 1 0 1052 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1269
timestamp 1524952243
transform 1 0 1116 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1296
timestamp 1524952243
transform 1 0 1012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1524952243
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1524952243
transform 1 0 1044 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1335
timestamp 1524952243
transform 1 0 980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1524952243
transform 1 0 1052 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1299
timestamp 1524952243
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1312
timestamp 1524952243
transform 1 0 1084 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1300
timestamp 1524952243
transform 1 0 1092 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1352
timestamp 1524952243
transform 1 0 1044 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1524952243
transform 1 0 1012 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1524952243
transform 1 0 1140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1524952243
transform 1 0 1148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1524952243
transform 1 0 1156 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1297
timestamp 1524952243
transform 1 0 1164 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1238
timestamp 1524952243
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1524952243
transform 1 0 1132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1524952243
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1524952243
transform 1 0 1164 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1353
timestamp 1524952243
transform 1 0 1124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1524952243
transform 1 0 1172 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1524952243
transform 1 0 1212 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1524952243
transform 1 0 1260 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1524952243
transform 1 0 1268 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1524952243
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1524952243
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1298
timestamp 1524952243
transform 1 0 1220 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1241
timestamp 1524952243
transform 1 0 1236 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1299
timestamp 1524952243
transform 1 0 1244 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1242
timestamp 1524952243
transform 1 0 1252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1524952243
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1524952243
transform 1 0 1188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1524952243
transform 1 0 1204 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1314
timestamp 1524952243
transform 1 0 1212 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1306
timestamp 1524952243
transform 1 0 1220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1524952243
transform 1 0 1228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1524952243
transform 1 0 1244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1524952243
transform 1 0 1268 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1354
timestamp 1524952243
transform 1 0 1188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1524952243
transform 1 0 1148 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1524952243
transform 1 0 1164 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1524952243
transform 1 0 1236 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1524952243
transform 1 0 1228 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1524952243
transform 1 0 1284 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1524952243
transform 1 0 1308 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1524952243
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1315
timestamp 1524952243
transform 1 0 1300 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1339
timestamp 1524952243
transform 1 0 1292 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_1356
timestamp 1524952243
transform 1 0 1284 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1524952243
transform 1 0 1332 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1524952243
transform 1 0 1356 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1524952243
transform 1 0 1348 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1311
timestamp 1524952243
transform 1 0 1340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1524952243
transform 1 0 1316 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1524952243
transform 1 0 1324 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1524952243
transform 1 0 1308 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_1357
timestamp 1524952243
transform 1 0 1324 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1524952243
transform 1 0 1348 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1524952243
transform 1 0 1396 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1524952243
transform 1 0 1388 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1524952243
transform 1 0 1388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1524952243
transform 1 0 1372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1524952243
transform 1 0 1348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1524952243
transform 1 0 1356 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1524952243
transform 1 0 1332 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_1358
timestamp 1524952243
transform 1 0 1348 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1524952243
transform 1 0 1460 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1524952243
transform 1 0 1468 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1524952243
transform 1 0 1452 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1245
timestamp 1524952243
transform 1 0 1436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1524952243
transform 1 0 1444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1524952243
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1524952243
transform 1 0 1468 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_1317
timestamp 1524952243
transform 1 0 1420 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1344
timestamp 1524952243
transform 1 0 1380 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1524952243
transform 1 0 1364 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_1373
timestamp 1524952243
transform 1 0 1340 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1524952243
transform 1 0 1316 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1524952243
transform 1 0 1380 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_1313
timestamp 1524952243
transform 1 0 1460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1318
timestamp 1524952243
transform 1 0 1468 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1524952243
transform 1 0 1508 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1524952243
transform 1 0 1492 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1524952243
transform 1 0 1524 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1524952243
transform 1 0 1556 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1524952243
transform 1 0 1620 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1524952243
transform 1 0 1628 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1524952243
transform 1 0 1596 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1249
timestamp 1524952243
transform 1 0 1492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1524952243
transform 1 0 1524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1524952243
transform 1 0 1532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1524952243
transform 1 0 1548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1524952243
transform 1 0 1556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1524952243
transform 1 0 1572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1524952243
transform 1 0 1588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1524952243
transform 1 0 1596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1524952243
transform 1 0 1476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1524952243
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1524952243
transform 1 0 1500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1524952243
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1524952243
transform 1 0 1524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1524952243
transform 1 0 1540 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1319
timestamp 1524952243
transform 1 0 1556 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1320
timestamp 1524952243
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1320
timestamp 1524952243
transform 1 0 1572 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1524952243
transform 1 0 1652 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1257
timestamp 1524952243
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1524952243
transform 1 0 1660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1524952243
transform 1 0 1580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1524952243
transform 1 0 1604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1336
timestamp 1524952243
transform 1 0 1492 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1524952243
transform 1 0 1524 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1524952243
transform 1 0 1556 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1524952243
transform 1 0 1500 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1524952243
transform 1 0 1540 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1524952243
transform 1 0 1628 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1323
timestamp 1524952243
transform 1 0 1636 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1322
timestamp 1524952243
transform 1 0 1652 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1524952243
transform 1 0 1684 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1524952243
transform 1 0 1684 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1524952243
transform 1 0 1692 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1524952243
transform 1 0 1756 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1524952243
transform 1 0 1804 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1524952243
transform 1 0 1740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1524952243
transform 1 0 1668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1524952243
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1524952243
transform 1 0 1692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1524952243
transform 1 0 1716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1524952243
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1361
timestamp 1524952243
transform 1 0 1596 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1524952243
transform 1 0 1660 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1524952243
transform 1 0 1676 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1524952243
transform 1 0 1580 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1524952243
transform 1 0 1604 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1524952243
transform 1 0 1588 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1524952243
transform 1 0 1716 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1524952243
transform 1 0 1796 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_1260
timestamp 1524952243
transform 1 0 1796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1524952243
transform 1 0 1772 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1323
timestamp 1524952243
transform 1 0 1780 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1524952243
transform 1 0 1796 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1330
timestamp 1524952243
transform 1 0 1804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1524952243
transform 1 0 1836 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1339
timestamp 1524952243
transform 1 0 1772 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1524952243
transform 1 0 1788 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1524952243
transform 1 0 1836 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1524952243
transform 1 0 1892 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1524952243
transform 1 0 1876 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1524952243
transform 1 0 2012 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1524952243
transform 1 0 1900 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1524952243
transform 1 0 1916 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1524952243
transform 1 0 1868 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1524952243
transform 1 0 1884 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1524952243
transform 1 0 1940 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1524952243
transform 1 0 1876 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_1261
timestamp 1524952243
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1524952243
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1524952243
transform 1 0 1940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1524952243
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1325
timestamp 1524952243
transform 1 0 1892 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_1333
timestamp 1524952243
transform 1 0 1916 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_1326
timestamp 1524952243
transform 1 0 1924 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1524952243
transform 1 0 1868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1524952243
transform 1 0 1916 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1524952243
transform 1 0 1908 0 1 905
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_20
timestamp 1524952243
transform 1 0 24 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_1387
timestamp 1524952243
transform 1 0 76 0 1 875
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_63
timestamp 1524952243
transform -1 0 168 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_56
timestamp 1524952243
transform -1 0 200 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1524952243
transform -1 0 232 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_85
timestamp 1524952243
transform 1 0 232 0 -1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_58
timestamp 1524952243
transform -1 0 280 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1524952243
transform -1 0 312 0 -1 970
box -8 -3 34 105
use NOR2X1  NOR2X1_31
timestamp 1524952243
transform 1 0 312 0 -1 970
box -8 -3 32 105
use INVX2  INVX2_86
timestamp 1524952243
transform 1 0 336 0 -1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_32
timestamp 1524952243
transform -1 0 392 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_87
timestamp 1524952243
transform 1 0 392 0 -1 970
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_64
timestamp 1524952243
transform 1 0 408 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_88
timestamp 1524952243
transform 1 0 504 0 -1 970
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_65
timestamp 1524952243
transform 1 0 520 0 -1 970
box -8 -3 104 105
use OAI22X1  OAI22X1_8
timestamp 1524952243
transform 1 0 616 0 -1 970
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_66
timestamp 1524952243
transform 1 0 656 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_89
timestamp 1524952243
transform 1 0 752 0 -1 970
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_67
timestamp 1524952243
transform 1 0 768 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_90
timestamp 1524952243
transform -1 0 880 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1524952243
transform 1 0 880 0 -1 970
box -9 -3 26 105
use M3_M2  M3_M2_1388
timestamp 1524952243
transform 1 0 932 0 1 875
box -3 -3 3 3
use OR2X1  OR2X1_4
timestamp 1524952243
transform 1 0 896 0 -1 970
box -8 -3 40 105
use OAI21X1  OAI21X1_60
timestamp 1524952243
transform 1 0 928 0 -1 970
box -8 -3 34 105
use NOR2X1  NOR2X1_32
timestamp 1524952243
transform -1 0 984 0 -1 970
box -8 -3 32 105
use XOR2X1  XOR2X1_21
timestamp 1524952243
transform -1 0 1040 0 -1 970
box -8 -3 64 105
use INVX2  INVX2_92
timestamp 1524952243
transform -1 0 1056 0 -1 970
box -9 -3 26 105
use XNOR2X1  XNOR2X1_17
timestamp 1524952243
transform 1 0 1056 0 -1 970
box -8 -3 64 105
use AND2X2  AND2X2_17
timestamp 1524952243
transform -1 0 1144 0 -1 970
box -8 -3 40 105
use AOI22X1  AOI22X1_33
timestamp 1524952243
transform -1 0 1184 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1524952243
transform 1 0 1184 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1524952243
transform 1 0 1224 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_1389
timestamp 1524952243
transform 1 0 1292 0 1 875
box -3 -3 3 3
use NOR2X1  NOR2X1_33
timestamp 1524952243
transform 1 0 1264 0 -1 970
box -8 -3 32 105
use NAND3X1  NAND3X1_18
timestamp 1524952243
transform -1 0 1320 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1524952243
transform -1 0 1352 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1524952243
transform -1 0 1384 0 -1 970
box -8 -3 40 105
use XNOR2X1  XNOR2X1_18
timestamp 1524952243
transform 1 0 1384 0 -1 970
box -8 -3 64 105
use AOI22X1  AOI22X1_36
timestamp 1524952243
transform -1 0 1480 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_1390
timestamp 1524952243
transform 1 0 1540 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_37
timestamp 1524952243
transform 1 0 1480 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1524952243
transform 1 0 1520 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1524952243
transform 1 0 1560 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_1391
timestamp 1524952243
transform 1 0 1660 0 1 875
box -3 -3 3 3
use XNOR2X1  XNOR2X1_19
timestamp 1524952243
transform 1 0 1600 0 -1 970
box -8 -3 64 105
use AND2X2  AND2X2_18
timestamp 1524952243
transform 1 0 1656 0 -1 970
box -8 -3 40 105
use XOR2X1  XOR2X1_22
timestamp 1524952243
transform 1 0 1688 0 -1 970
box -8 -3 64 105
use M3_M2  M3_M2_1392
timestamp 1524952243
transform 1 0 1756 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1524952243
transform 1 0 1772 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_23
timestamp 1524952243
transform 1 0 1744 0 -1 970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_20
timestamp 1524952243
transform 1 0 1800 0 -1 970
box -8 -3 64 105
use AND2X2  AND2X2_19
timestamp 1524952243
transform -1 0 1888 0 -1 970
box -8 -3 40 105
use M3_M2  M3_M2_1394
timestamp 1524952243
transform 1 0 1908 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_24
timestamp 1524952243
transform 1 0 1888 0 -1 970
box -8 -3 64 105
use top_module_VIA0  top_module_VIA0_21
timestamp 1524952243
transform 1 0 1994 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_1403
timestamp 1524952243
transform 1 0 68 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1524952243
transform 1 0 204 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_1350
timestamp 1524952243
transform 1 0 172 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1524952243
transform 1 0 68 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1474
timestamp 1524952243
transform 1 0 76 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1362
timestamp 1524952243
transform 1 0 124 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1447
timestamp 1524952243
transform 1 0 196 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1524952243
transform 1 0 204 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1524952243
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1524952243
transform 1 0 196 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1475
timestamp 1524952243
transform 1 0 204 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1524952243
transform 1 0 228 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1524952243
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1524952243
transform 1 0 156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1524952243
transform 1 0 172 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1496
timestamp 1524952243
transform 1 0 180 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1524952243
transform 1 0 196 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1437
timestamp 1524952243
transform 1 0 204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1524952243
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1524952243
transform 1 0 236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1524952243
transform 1 0 236 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_1540
timestamp 1524952243
transform 1 0 228 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1524952243
transform 1 0 252 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1366
timestamp 1524952243
transform 1 0 252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1524952243
transform 1 0 252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1524952243
transform 1 0 260 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_1541
timestamp 1524952243
transform 1 0 252 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1352
timestamp 1524952243
transform 1 0 284 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_1448
timestamp 1524952243
transform 1 0 300 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1353
timestamp 1524952243
transform 1 0 308 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1524952243
transform 1 0 276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1524952243
transform 1 0 292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1524952243
transform 1 0 300 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1498
timestamp 1524952243
transform 1 0 276 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1441
timestamp 1524952243
transform 1 0 300 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1516
timestamp 1524952243
transform 1 0 300 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1524952243
transform 1 0 324 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1524952243
transform 1 0 332 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1524952243
transform 1 0 396 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1524952243
transform 1 0 380 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1524952243
transform 1 0 388 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1370
timestamp 1524952243
transform 1 0 340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1524952243
transform 1 0 348 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1524952243
transform 1 0 356 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1524952243
transform 1 0 420 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1372
timestamp 1524952243
transform 1 0 364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1524952243
transform 1 0 380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1524952243
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1524952243
transform 1 0 404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1524952243
transform 1 0 324 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1499
timestamp 1524952243
transform 1 0 340 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1443
timestamp 1524952243
transform 1 0 356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1500
timestamp 1524952243
transform 1 0 364 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1524952243
transform 1 0 412 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1376
timestamp 1524952243
transform 1 0 420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1524952243
transform 1 0 428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1524952243
transform 1 0 388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1524952243
transform 1 0 396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1524952243
transform 1 0 412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1524952243
transform 1 0 420 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1524952243
transform 1 0 324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1524952243
transform 1 0 388 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1524952243
transform 1 0 508 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1524952243
transform 1 0 460 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1524952243
transform 1 0 452 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1524952243
transform 1 0 492 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1524952243
transform 1 0 436 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1448
timestamp 1524952243
transform 1 0 444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1524952243
transform 1 0 452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1524952243
transform 1 0 492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1524952243
transform 1 0 556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1524952243
transform 1 0 468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1524952243
transform 1 0 556 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1543
timestamp 1524952243
transform 1 0 556 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1524952243
transform 1 0 580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1524952243
transform 1 0 596 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1524952243
transform 1 0 572 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1381
timestamp 1524952243
transform 1 0 572 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1502
timestamp 1524952243
transform 1 0 564 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1451
timestamp 1524952243
transform 1 0 572 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1518
timestamp 1524952243
transform 1 0 564 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1382
timestamp 1524952243
transform 1 0 580 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1478
timestamp 1524952243
transform 1 0 588 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1383
timestamp 1524952243
transform 1 0 596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1524952243
transform 1 0 588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1503
timestamp 1524952243
transform 1 0 596 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1524952243
transform 1 0 628 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1524952243
transform 1 0 636 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1524952243
transform 1 0 708 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1524952243
transform 1 0 676 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1385
timestamp 1524952243
transform 1 0 644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1524952243
transform 1 0 660 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1480
timestamp 1524952243
transform 1 0 668 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1524952243
transform 1 0 724 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1387
timestamp 1524952243
transform 1 0 684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1524952243
transform 1 0 700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1524952243
transform 1 0 636 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1504
timestamp 1524952243
transform 1 0 644 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1524952243
transform 1 0 708 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1389
timestamp 1524952243
transform 1 0 716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1524952243
transform 1 0 772 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1482
timestamp 1524952243
transform 1 0 796 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1454
timestamp 1524952243
transform 1 0 652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1524952243
transform 1 0 668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1524952243
transform 1 0 676 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1519
timestamp 1524952243
transform 1 0 612 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1524952243
transform 1 0 628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1524952243
transform 1 0 684 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1524952243
transform 1 0 940 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1524952243
transform 1 0 932 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1524952243
transform 1 0 940 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1524952243
transform 1 0 876 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1524952243
transform 1 0 900 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1524952243
transform 1 0 948 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1391
timestamp 1524952243
transform 1 0 820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1524952243
transform 1 0 836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1524952243
transform 1 0 844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1524952243
transform 1 0 692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1524952243
transform 1 0 708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1524952243
transform 1 0 796 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1524952243
transform 1 0 812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1524952243
transform 1 0 828 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1521
timestamp 1524952243
transform 1 0 668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1524952243
transform 1 0 684 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1524952243
transform 1 0 724 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1524952243
transform 1 0 772 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1524952243
transform 1 0 836 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1524952243
transform 1 0 860 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1524952243
transform 1 0 892 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1394
timestamp 1524952243
transform 1 0 900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1524952243
transform 1 0 940 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1485
timestamp 1524952243
transform 1 0 948 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1524952243
transform 1 0 1004 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1524952243
transform 1 0 988 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1524952243
transform 1 0 1044 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1524952243
transform 1 0 1044 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1524952243
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1524952243
transform 1 0 972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1524952243
transform 1 0 988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1524952243
transform 1 0 1004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1524952243
transform 1 0 1036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1524952243
transform 1 0 860 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1507
timestamp 1524952243
transform 1 0 884 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1463
timestamp 1524952243
transform 1 0 948 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1525
timestamp 1524952243
transform 1 0 828 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1524952243
transform 1 0 844 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1524952243
transform 1 0 876 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1524952243
transform 1 0 900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1524952243
transform 1 0 708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1524952243
transform 1 0 772 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1524952243
transform 1 0 812 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1524952243
transform 1 0 908 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1524952243
transform 1 0 956 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1524952243
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1524952243
transform 1 0 980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1524952243
transform 1 0 988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1524952243
transform 1 0 1036 0 1 807
box -2 -2 2 2
use M3_M2  M3_M2_1529
timestamp 1524952243
transform 1 0 964 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1524952243
transform 1 0 980 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1524952243
transform 1 0 1028 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1524952243
transform 1 0 1068 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1524952243
transform 1 0 1060 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1524952243
transform 1 0 1108 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1524952243
transform 1 0 1092 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1401
timestamp 1524952243
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1524952243
transform 1 0 1060 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1524952243
transform 1 0 1244 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1524952243
transform 1 0 1124 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1348
timestamp 1524952243
transform 1 0 1140 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_1436
timestamp 1524952243
transform 1 0 1148 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1524952243
transform 1 0 1164 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1524952243
transform 1 0 1180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1524952243
transform 1 0 1212 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1524952243
transform 1 0 1108 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1524952243
transform 1 0 1124 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1524952243
transform 1 0 1100 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1467
timestamp 1524952243
transform 1 0 1076 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1510
timestamp 1524952243
transform 1 0 1084 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1434
timestamp 1524952243
transform 1 0 1100 0 1 807
box -2 -2 2 2
use M3_M2  M3_M2_1530
timestamp 1524952243
transform 1 0 1076 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1524952243
transform 1 0 1140 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1357
timestamp 1524952243
transform 1 0 1148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1524952243
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1524952243
transform 1 0 1148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1524952243
transform 1 0 1124 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1511
timestamp 1524952243
transform 1 0 1132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1524952243
transform 1 0 1300 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1524952243
transform 1 0 1276 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1524952243
transform 1 0 1372 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1524952243
transform 1 0 1308 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1524952243
transform 1 0 1332 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1524952243
transform 1 0 1364 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1524952243
transform 1 0 1284 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1524952243
transform 1 0 1220 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1524952243
transform 1 0 1244 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1524952243
transform 1 0 1276 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1524952243
transform 1 0 1316 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1404
timestamp 1524952243
transform 1 0 1196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1524952243
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1524952243
transform 1 0 1244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1524952243
transform 1 0 1276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1524952243
transform 1 0 1292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1524952243
transform 1 0 1308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1524952243
transform 1 0 1316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1524952243
transform 1 0 1164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1524952243
transform 1 0 1220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1524952243
transform 1 0 1276 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1512
timestamp 1524952243
transform 1 0 1292 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1524952243
transform 1 0 1332 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1524952243
transform 1 0 1524 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1524952243
transform 1 0 1476 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1524952243
transform 1 0 1444 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1524952243
transform 1 0 1436 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1524952243
transform 1 0 1476 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1524952243
transform 1 0 1396 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1524952243
transform 1 0 1420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1524952243
transform 1 0 1460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1524952243
transform 1 0 1532 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1524952243
transform 1 0 1564 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_1411
timestamp 1524952243
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1524952243
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1524952243
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1524952243
transform 1 0 1420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1524952243
transform 1 0 1444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1524952243
transform 1 0 1476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1524952243
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1524952243
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1524952243
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1524952243
transform 1 0 1284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1524952243
transform 1 0 1308 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1474
timestamp 1524952243
transform 1 0 1372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1531
timestamp 1524952243
transform 1 0 1364 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1475
timestamp 1524952243
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1489
timestamp 1524952243
transform 1 0 1508 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1524952243
transform 1 0 1476 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1476
timestamp 1524952243
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1552
timestamp 1524952243
transform 1 0 1372 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1524952243
transform 1 0 1388 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1524952243
transform 1 0 1420 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1524952243
transform 1 0 1444 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1524952243
transform 1 0 1572 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1418
timestamp 1524952243
transform 1 0 1564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1524952243
transform 1 0 1572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1524952243
transform 1 0 1532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1524952243
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1467
timestamp 1524952243
transform 1 0 1644 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1524952243
transform 1 0 1620 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1524952243
transform 1 0 1716 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1524952243
transform 1 0 1748 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1524952243
transform 1 0 1724 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1524952243
transform 1 0 1772 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1524952243
transform 1 0 1692 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1524952243
transform 1 0 1740 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1524952243
transform 1 0 1764 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1420
timestamp 1524952243
transform 1 0 1644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1524952243
transform 1 0 1652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1524952243
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1524952243
transform 1 0 1692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1524952243
transform 1 0 1588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1514
timestamp 1524952243
transform 1 0 1596 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1524952243
transform 1 0 1596 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1524952243
transform 1 0 1492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1524952243
transform 1 0 1524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1524952243
transform 1 0 1540 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1524952243
transform 1 0 1572 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1480
timestamp 1524952243
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1524952243
transform 1 0 1652 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1515
timestamp 1524952243
transform 1 0 1668 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1524952243
transform 1 0 1716 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1524952243
transform 1 0 1724 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1492
timestamp 1524952243
transform 1 0 1740 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1524952243
transform 1 0 1804 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1524952243
transform 1 0 1796 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1524952243
transform 1 0 1820 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1524952243
transform 1 0 1852 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1524952243
transform 1 0 1852 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1524952243
transform 1 0 1876 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_1349
timestamp 1524952243
transform 1 0 1852 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_1446
timestamp 1524952243
transform 1 0 1860 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1358
timestamp 1524952243
transform 1 0 1836 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1524952243
transform 1 0 1844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1524952243
transform 1 0 1748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1524952243
transform 1 0 1764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1524952243
transform 1 0 1676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1524952243
transform 1 0 1684 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1533
timestamp 1524952243
transform 1 0 1660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1524952243
transform 1 0 1684 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1524952243
transform 1 0 1780 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1427
timestamp 1524952243
transform 1 0 1788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1524952243
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1524952243
transform 1 0 1748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1524952243
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1524952243
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1524952243
transform 1 0 1780 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1535
timestamp 1524952243
transform 1 0 1748 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1524952243
transform 1 0 1708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1524952243
transform 1 0 1780 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1524952243
transform 1 0 1780 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1429
timestamp 1524952243
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1524952243
transform 1 0 1812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1524952243
transform 1 0 1820 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1537
timestamp 1524952243
transform 1 0 1812 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1524952243
transform 1 0 1828 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1360
timestamp 1524952243
transform 1 0 1868 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_1494
timestamp 1524952243
transform 1 0 1852 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1430
timestamp 1524952243
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1524952243
transform 1 0 1876 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_1473
timestamp 1524952243
transform 1 0 1908 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1524952243
transform 1 0 1924 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1432
timestamp 1524952243
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1524952243
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1524952243
transform 1 0 1892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1524952243
transform 1 0 1940 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_1539
timestamp 1524952243
transform 1 0 1860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1524952243
transform 1 0 1844 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1524952243
transform 1 0 1932 0 1 785
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_22
timestamp 1524952243
transform 1 0 48 0 1 770
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_68
timestamp 1524952243
transform -1 0 168 0 1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_61
timestamp 1524952243
transform -1 0 200 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_1564
timestamp 1524952243
transform 1 0 212 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1524952243
transform 1 0 236 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_62
timestamp 1524952243
transform -1 0 232 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_1566
timestamp 1524952243
transform 1 0 260 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_34
timestamp 1524952243
transform 1 0 232 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_1567
timestamp 1524952243
transform 1 0 276 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_35
timestamp 1524952243
transform 1 0 256 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1524952243
transform -1 0 304 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1524952243
transform -1 0 328 0 1 770
box -8 -3 32 105
use INVX2  INVX2_93
timestamp 1524952243
transform 1 0 328 0 1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_40
timestamp 1524952243
transform -1 0 384 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_1568
timestamp 1524952243
transform 1 0 428 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_41
timestamp 1524952243
transform -1 0 424 0 1 770
box -8 -3 46 105
use INVX2  INVX2_94
timestamp 1524952243
transform 1 0 424 0 1 770
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1524952243
transform 1 0 440 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_1569
timestamp 1524952243
transform 1 0 516 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1524952243
transform 1 0 556 0 1 775
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_69
timestamp 1524952243
transform 1 0 456 0 1 770
box -8 -3 104 105
use INVX2  INVX2_96
timestamp 1524952243
transform 1 0 552 0 1 770
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1524952243
transform 1 0 568 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_1571
timestamp 1524952243
transform 1 0 604 0 1 775
box -3 -3 3 3
use AND2X2  AND2X2_20
timestamp 1524952243
transform 1 0 584 0 1 770
box -8 -3 40 105
use INVX2  INVX2_98
timestamp 1524952243
transform 1 0 616 0 1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_9
timestamp 1524952243
transform 1 0 632 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1524952243
transform 1 0 672 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_1572
timestamp 1524952243
transform 1 0 756 0 1 775
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_70
timestamp 1524952243
transform -1 0 808 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_1573
timestamp 1524952243
transform 1 0 828 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_11
timestamp 1524952243
transform -1 0 848 0 1 770
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_71
timestamp 1524952243
transform 1 0 848 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_1574
timestamp 1524952243
transform 1 0 972 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_12
timestamp 1524952243
transform 1 0 944 0 1 770
box -8 -3 46 105
use XNOR2X1  XNOR2X1_21
timestamp 1524952243
transform -1 0 1040 0 1 770
box -8 -3 64 105
use OAI21X1  OAI21X1_63
timestamp 1524952243
transform -1 0 1072 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1524952243
transform 1 0 1072 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_1575
timestamp 1524952243
transform 1 0 1124 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_34
timestamp 1524952243
transform -1 0 1128 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_1576
timestamp 1524952243
transform 1 0 1148 0 1 775
box -3 -3 3 3
use NAND3X1  NAND3X1_21
timestamp 1524952243
transform -1 0 1160 0 1 770
box -8 -3 40 105
use M3_M2  M3_M2_1577
timestamp 1524952243
transform 1 0 1220 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_25
timestamp 1524952243
transform 1 0 1160 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_1578
timestamp 1524952243
transform 1 0 1276 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_26
timestamp 1524952243
transform 1 0 1216 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_1579
timestamp 1524952243
transform 1 0 1300 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1524952243
transform 1 0 1316 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_42
timestamp 1524952243
transform -1 0 1312 0 1 770
box -8 -3 46 105
use XNOR2X1  XNOR2X1_22
timestamp 1524952243
transform -1 0 1368 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_27
timestamp 1524952243
transform 1 0 1368 0 1 770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_23
timestamp 1524952243
transform -1 0 1480 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_28
timestamp 1524952243
transform -1 0 1536 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_29
timestamp 1524952243
transform 1 0 1536 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_1581
timestamp 1524952243
transform 1 0 1644 0 1 775
box -3 -3 3 3
use XNOR2X1  XNOR2X1_24
timestamp 1524952243
transform 1 0 1592 0 1 770
box -8 -3 64 105
use AOI22X1  AOI22X1_43
timestamp 1524952243
transform -1 0 1688 0 1 770
box -8 -3 46 105
use XOR2X1  XOR2X1_30
timestamp 1524952243
transform 1 0 1688 0 1 770
box -8 -3 64 105
use AOI22X1  AOI22X1_44
timestamp 1524952243
transform -1 0 1784 0 1 770
box -8 -3 46 105
use OAI21X1  OAI21X1_65
timestamp 1524952243
transform 1 0 1784 0 1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_35
timestamp 1524952243
transform 1 0 1816 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_1582
timestamp 1524952243
transform 1 0 1852 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1524952243
transform 1 0 1868 0 1 775
box -3 -3 3 3
use NAND3X1  NAND3X1_22
timestamp 1524952243
transform -1 0 1872 0 1 770
box -8 -3 40 105
use M3_M2  M3_M2_1584
timestamp 1524952243
transform 1 0 1892 0 1 775
box -3 -3 3 3
use INVX2  INVX2_99
timestamp 1524952243
transform -1 0 1888 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_1585
timestamp 1524952243
transform 1 0 1908 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1524952243
transform 1 0 1940 0 1 775
box -3 -3 3 3
use XNOR2X1  XNOR2X1_25
timestamp 1524952243
transform 1 0 1888 0 1 770
box -8 -3 64 105
use top_module_VIA0  top_module_VIA0_23
timestamp 1524952243
transform 1 0 1970 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_1609
timestamp 1524952243
transform 1 0 68 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1552
timestamp 1524952243
transform 1 0 76 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1748
timestamp 1524952243
transform 1 0 68 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1524952243
transform 1 0 148 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1524952243
transform 1 0 172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1498
timestamp 1524952243
transform 1 0 172 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1665
timestamp 1524952243
transform 1 0 132 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1499
timestamp 1524952243
transform 1 0 220 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1649
timestamp 1524952243
transform 1 0 228 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1524952243
transform 1 0 268 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1524952243
transform 1 0 268 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1500
timestamp 1524952243
transform 1 0 244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1524952243
transform 1 0 148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1524952243
transform 1 0 188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1694
timestamp 1524952243
transform 1 0 140 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1524952243
transform 1 0 172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1524952243
transform 1 0 196 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1555
timestamp 1524952243
transform 1 0 204 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1524952243
transform 1 0 220 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1524952243
transform 1 0 252 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1501
timestamp 1524952243
transform 1 0 268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1524952243
transform 1 0 228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1524952243
transform 1 0 244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1524952243
transform 1 0 252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1524952243
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1524952243
transform 1 0 188 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1524952243
transform 1 0 220 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1749
timestamp 1524952243
transform 1 0 220 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_1625
timestamp 1524952243
transform 1 0 268 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1524952243
transform 1 0 284 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1668
timestamp 1524952243
transform 1 0 284 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1524952243
transform 1 0 308 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1524952243
transform 1 0 316 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1560
timestamp 1524952243
transform 1 0 300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1524952243
transform 1 0 284 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1721
timestamp 1524952243
transform 1 0 284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1524952243
transform 1 0 308 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1561
timestamp 1524952243
transform 1 0 316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1524952243
transform 1 0 308 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1629
timestamp 1524952243
transform 1 0 340 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1503
timestamp 1524952243
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1524952243
transform 1 0 356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1524952243
transform 1 0 364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1524952243
transform 1 0 324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1524952243
transform 1 0 332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1524952243
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1524952243
transform 1 0 364 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1670
timestamp 1524952243
transform 1 0 372 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1524952243
transform 1 0 436 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1524952243
transform 1 0 404 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1506
timestamp 1524952243
transform 1 0 468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1524952243
transform 1 0 380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1524952243
transform 1 0 388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1524952243
transform 1 0 428 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1722
timestamp 1524952243
transform 1 0 356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1524952243
transform 1 0 380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1524952243
transform 1 0 428 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1524952243
transform 1 0 388 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1524952243
transform 1 0 364 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1524952243
transform 1 0 396 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1524952243
transform 1 0 444 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1524952243
transform 1 0 340 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1524952243
transform 1 0 524 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1524952243
transform 1 0 548 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1524952243
transform 1 0 540 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1507
timestamp 1524952243
transform 1 0 492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1524952243
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1524952243
transform 1 0 572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1524952243
transform 1 0 580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1698
timestamp 1524952243
transform 1 0 580 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1524952243
transform 1 0 524 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1524952243
transform 1 0 588 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1524952243
transform 1 0 620 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1524952243
transform 1 0 668 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1524952243
transform 1 0 604 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1524952243
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1524952243
transform 1 0 596 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1737
timestamp 1524952243
transform 1 0 596 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_1508
timestamp 1524952243
transform 1 0 620 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1653
timestamp 1524952243
transform 1 0 660 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1524952243
transform 1 0 604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1524952243
transform 1 0 652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1524952243
transform 1 0 700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1524952243
transform 1 0 708 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1699
timestamp 1524952243
transform 1 0 644 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1524952243
transform 1 0 700 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1524952243
transform 1 0 716 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_1509
timestamp 1524952243
transform 1 0 716 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1671
timestamp 1524952243
transform 1 0 716 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1578
timestamp 1524952243
transform 1 0 724 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1725
timestamp 1524952243
transform 1 0 724 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1524952243
transform 1 0 732 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1524952243
transform 1 0 740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1524952243
transform 1 0 756 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1524952243
transform 1 0 732 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1524952243
transform 1 0 876 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1524952243
transform 1 0 812 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1524952243
transform 1 0 868 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1524952243
transform 1 0 916 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1510
timestamp 1524952243
transform 1 0 740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1524952243
transform 1 0 756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1524952243
transform 1 0 772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1524952243
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1524952243
transform 1 0 876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1524952243
transform 1 0 892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1524952243
transform 1 0 908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1524952243
transform 1 0 916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1524952243
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1524952243
transform 1 0 740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1672
timestamp 1524952243
transform 1 0 748 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1581
timestamp 1524952243
transform 1 0 764 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1673
timestamp 1524952243
transform 1 0 772 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1524952243
transform 1 0 788 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1582
timestamp 1524952243
transform 1 0 812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1524952243
transform 1 0 868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1524952243
transform 1 0 884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1524952243
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1524952243
transform 1 0 916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1700
timestamp 1524952243
transform 1 0 740 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1524952243
transform 1 0 764 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1524952243
transform 1 0 788 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1524952243
transform 1 0 828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1524952243
transform 1 0 788 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1524952243
transform 1 0 916 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1524952243
transform 1 0 1020 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1524952243
transform 1 0 1060 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1524952243
transform 1 0 996 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1524952243
transform 1 0 988 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1518
timestamp 1524952243
transform 1 0 988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1524952243
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1524952243
transform 1 0 1020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1524952243
transform 1 0 948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1524952243
transform 1 0 980 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1521
timestamp 1524952243
transform 1 0 1076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1524952243
transform 1 0 988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1524952243
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1524952243
transform 1 0 1028 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1703
timestamp 1524952243
transform 1 0 948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1524952243
transform 1 0 924 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1524952243
transform 1 0 956 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1524952243
transform 1 0 996 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1524952243
transform 1 0 1012 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1524952243
transform 1 0 1052 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1524952243
transform 1 0 1140 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_1591
timestamp 1524952243
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1524952243
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1705
timestamp 1524952243
transform 1 0 1060 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1524952243
transform 1 0 1108 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1593
timestamp 1524952243
transform 1 0 1116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1739
timestamp 1524952243
transform 1 0 1052 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1524952243
transform 1 0 1076 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1524952243
transform 1 0 1068 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1524952243
transform 1 0 1172 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1524952243
transform 1 0 1212 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1524952243
transform 1 0 1164 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1524952243
transform 1 0 1148 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1524952243
transform 1 0 1164 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1524952243
transform 1 0 1156 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1522
timestamp 1524952243
transform 1 0 1164 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1656
timestamp 1524952243
transform 1 0 1172 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1524952243
transform 1 0 1220 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1524952243
transform 1 0 1268 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1523
timestamp 1524952243
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1524952243
transform 1 0 1236 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1657
timestamp 1524952243
transform 1 0 1244 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1594
timestamp 1524952243
transform 1 0 1156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1524952243
transform 1 0 1172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1524952243
transform 1 0 1196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1524952243
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1706
timestamp 1524952243
transform 1 0 1132 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1524952243
transform 1 0 1196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1524952243
transform 1 0 1236 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1495
timestamp 1524952243
transform 1 0 1300 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1524952243
transform 1 0 1332 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_1658
timestamp 1524952243
transform 1 0 1292 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1524952243
transform 1 0 1308 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1525
timestamp 1524952243
transform 1 0 1316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1524952243
transform 1 0 1324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1524952243
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1524952243
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1524952243
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1708
timestamp 1524952243
transform 1 0 1276 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1524952243
transform 1 0 1260 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1524952243
transform 1 0 1316 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1524952243
transform 1 0 1348 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1524952243
transform 1 0 1348 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1524952243
transform 1 0 1396 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1524952243
transform 1 0 1364 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1524952243
transform 1 0 1428 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1527
timestamp 1524952243
transform 1 0 1348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1524952243
transform 1 0 1380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1524952243
transform 1 0 1388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1524952243
transform 1 0 1396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1524952243
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1680
timestamp 1524952243
transform 1 0 1340 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1602
timestamp 1524952243
transform 1 0 1348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1524952243
transform 1 0 1356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1524952243
transform 1 0 1372 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1709
timestamp 1524952243
transform 1 0 1308 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1524952243
transform 1 0 1332 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1524952243
transform 1 0 1324 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1524952243
transform 1 0 1380 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1524952243
transform 1 0 1372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1524952243
transform 1 0 1476 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1524952243
transform 1 0 1492 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1524952243
transform 1 0 1484 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1524952243
transform 1 0 1452 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1524952243
transform 1 0 1444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1524952243
transform 1 0 1452 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1618
timestamp 1524952243
transform 1 0 1516 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1524952243
transform 1 0 1540 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1524952243
transform 1 0 1524 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1524952243
transform 1 0 1500 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1660
timestamp 1524952243
transform 1 0 1508 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1534
timestamp 1524952243
transform 1 0 1516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1524952243
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1524952243
transform 1 0 1532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1524952243
transform 1 0 1444 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1682
timestamp 1524952243
transform 1 0 1452 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1524952243
transform 1 0 1476 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1606
timestamp 1524952243
transform 1 0 1508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1524952243
transform 1 0 1524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1712
timestamp 1524952243
transform 1 0 1444 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1524952243
transform 1 0 1508 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1524952243
transform 1 0 1532 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1524952243
transform 1 0 1556 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1537
timestamp 1524952243
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1661
timestamp 1524952243
transform 1 0 1580 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1538
timestamp 1524952243
transform 1 0 1596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1524952243
transform 1 0 1548 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1685
timestamp 1524952243
transform 1 0 1564 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1628
timestamp 1524952243
transform 1 0 1532 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1729
timestamp 1524952243
transform 1 0 1516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1524952243
transform 1 0 1548 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1524952243
transform 1 0 1620 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1539
timestamp 1524952243
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1686
timestamp 1524952243
transform 1 0 1604 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1609
timestamp 1524952243
transform 1 0 1612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1524952243
transform 1 0 1620 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1687
timestamp 1524952243
transform 1 0 1628 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1629
timestamp 1524952243
transform 1 0 1564 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1524952243
transform 1 0 1588 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1524952243
transform 1 0 1596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1524952243
transform 1 0 1572 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_1730
timestamp 1524952243
transform 1 0 1580 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1524952243
transform 1 0 1572 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1524952243
transform 1 0 1628 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1604
timestamp 1524952243
transform 1 0 1676 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1524952243
transform 1 0 1668 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1540
timestamp 1524952243
transform 1 0 1644 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1605
timestamp 1524952243
transform 1 0 1740 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1524952243
transform 1 0 1748 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1524952243
transform 1 0 1700 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1541
timestamp 1524952243
transform 1 0 1708 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1688
timestamp 1524952243
transform 1 0 1644 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1524952243
transform 1 0 1676 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1689
timestamp 1524952243
transform 1 0 1684 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1524952243
transform 1 0 1796 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1524952243
transform 1 0 1828 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1524952243
transform 1 0 1796 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1524952243
transform 1 0 1812 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1542
timestamp 1524952243
transform 1 0 1764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1524952243
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1524952243
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1524952243
transform 1 0 1644 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1731
timestamp 1524952243
transform 1 0 1660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1524952243
transform 1 0 1732 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1543
timestamp 1524952243
transform 1 0 1812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1524952243
transform 1 0 1820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1524952243
transform 1 0 1740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1524952243
transform 1 0 1756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1524952243
transform 1 0 1788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1715
timestamp 1524952243
transform 1 0 1740 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1524952243
transform 1 0 1732 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1524952243
transform 1 0 1668 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1524952243
transform 1 0 1708 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1524952243
transform 1 0 1796 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1524952243
transform 1 0 1812 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1524952243
transform 1 0 1876 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1524952243
transform 1 0 1860 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1524952243
transform 1 0 1892 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1497
timestamp 1524952243
transform 1 0 1884 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1524952243
transform 1 0 1844 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1524952243
transform 1 0 1852 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1546
timestamp 1524952243
transform 1 0 1860 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_1664
timestamp 1524952243
transform 1 0 1884 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1524952243
transform 1 0 1900 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1524952243
transform 1 0 1924 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1547
timestamp 1524952243
transform 1 0 1892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1524952243
transform 1 0 1900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1524952243
transform 1 0 1916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1524952243
transform 1 0 1932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1524952243
transform 1 0 2012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1524952243
transform 1 0 1828 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1716
timestamp 1524952243
transform 1 0 1788 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1524952243
transform 1 0 1780 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1524952243
transform 1 0 1756 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1524952243
transform 1 0 1828 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1618
timestamp 1524952243
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1524952243
transform 1 0 1876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1524952243
transform 1 0 1844 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_1745
timestamp 1524952243
transform 1 0 1836 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1524952243
transform 1 0 1860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1524952243
transform 1 0 1876 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1524952243
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1524952243
transform 1 0 1924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1524952243
transform 1 0 1948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1693
timestamp 1524952243
transform 1 0 2012 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1524952243
transform 1 0 1932 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1524952243
transform 1 0 1916 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1524952243
transform 1 0 1948 0 1 695
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_24
timestamp 1524952243
transform 1 0 24 0 1 670
box -10 -3 10 3
use FILL  FILL_15
timestamp 1524952243
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_16
timestamp 1524952243
transform 1 0 80 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_1757
timestamp 1524952243
transform 1 0 108 0 1 675
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_72
timestamp 1524952243
transform -1 0 184 0 -1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_66
timestamp 1524952243
transform -1 0 216 0 -1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_36
timestamp 1524952243
transform -1 0 240 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1524952243
transform 1 0 240 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1524952243
transform 1 0 264 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1524952243
transform 1 0 288 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_100
timestamp 1524952243
transform 1 0 312 0 -1 770
box -9 -3 26 105
use M3_M2  M3_M2_1758
timestamp 1524952243
transform 1 0 348 0 1 675
box -3 -3 3 3
use AOI22X1  AOI22X1_45
timestamp 1524952243
transform -1 0 368 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_101
timestamp 1524952243
transform 1 0 368 0 -1 770
box -9 -3 26 105
use M3_M2  M3_M2_1759
timestamp 1524952243
transform 1 0 428 0 1 675
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_73
timestamp 1524952243
transform -1 0 480 0 -1 770
box -8 -3 104 105
use M3_M2  M3_M2_1760
timestamp 1524952243
transform 1 0 564 0 1 675
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_74
timestamp 1524952243
transform 1 0 480 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_102
timestamp 1524952243
transform 1 0 576 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1524952243
transform 1 0 592 0 -1 770
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_75
timestamp 1524952243
transform 1 0 608 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_104
timestamp 1524952243
transform -1 0 720 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1524952243
transform 1 0 720 0 -1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_13
timestamp 1524952243
transform 1 0 736 0 -1 770
box -8 -3 46 105
use DFFPOSX1  DFFPOSX1_76
timestamp 1524952243
transform 1 0 776 0 -1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_14
timestamp 1524952243
transform 1 0 872 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_106
timestamp 1524952243
transform 1 0 912 0 -1 770
box -9 -3 26 105
use XNOR2X1  XNOR2X1_26
timestamp 1524952243
transform -1 0 984 0 -1 770
box -8 -3 64 105
use AOI22X1  AOI22X1_46
timestamp 1524952243
transform -1 0 1024 0 -1 770
box -8 -3 46 105
use XNOR2X1  XNOR2X1_27
timestamp 1524952243
transform 1 0 1024 0 -1 770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_28
timestamp 1524952243
transform 1 0 1080 0 -1 770
box -8 -3 64 105
use AND2X2  AND2X2_21
timestamp 1524952243
transform -1 0 1168 0 -1 770
box -8 -3 40 105
use XOR2X1  XOR2X1_31
timestamp 1524952243
transform 1 0 1168 0 -1 770
box -8 -3 64 105
use INVX2  INVX2_107
timestamp 1524952243
transform -1 0 1240 0 -1 770
box -9 -3 26 105
use XOR2X1  XOR2X1_32
timestamp 1524952243
transform 1 0 1240 0 -1 770
box -8 -3 64 105
use AOI21X1  AOI21X1_8
timestamp 1524952243
transform -1 0 1328 0 -1 770
box -7 -3 39 105
use M3_M2  M3_M2_1761
timestamp 1524952243
transform 1 0 1356 0 1 675
box -3 -3 3 3
use NOR2X1  NOR2X1_36
timestamp 1524952243
transform 1 0 1328 0 -1 770
box -8 -3 32 105
use M3_M2  M3_M2_1762
timestamp 1524952243
transform 1 0 1388 0 1 675
box -3 -3 3 3
use AOI22X1  AOI22X1_47
timestamp 1524952243
transform 1 0 1352 0 -1 770
box -8 -3 46 105
use XNOR2X1  XNOR2X1_29
timestamp 1524952243
transform -1 0 1448 0 -1 770
box -8 -3 64 105
use M3_M2  M3_M2_1763
timestamp 1524952243
transform 1 0 1476 0 1 675
box -3 -3 3 3
use XNOR2X1  XNOR2X1_30
timestamp 1524952243
transform 1 0 1448 0 -1 770
box -8 -3 64 105
use NOR2X1  NOR2X1_37
timestamp 1524952243
transform 1 0 1504 0 -1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_67
timestamp 1524952243
transform -1 0 1560 0 -1 770
box -8 -3 34 105
use NAND3X1  NAND3X1_23
timestamp 1524952243
transform -1 0 1592 0 -1 770
box -8 -3 40 105
use OAI21X1  OAI21X1_68
timestamp 1524952243
transform -1 0 1624 0 -1 770
box -8 -3 34 105
use M3_M2  M3_M2_1764
timestamp 1524952243
transform 1 0 1644 0 1 675
box -3 -3 3 3
use NAND2X1  NAND2X1_40
timestamp 1524952243
transform -1 0 1648 0 -1 770
box -8 -3 32 105
use M3_M2  M3_M2_1765
timestamp 1524952243
transform 1 0 1692 0 1 675
box -3 -3 3 3
use XOR2X1  XOR2X1_33
timestamp 1524952243
transform 1 0 1648 0 -1 770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_31
timestamp 1524952243
transform 1 0 1704 0 -1 770
box -8 -3 64 105
use M3_M2  M3_M2_1766
timestamp 1524952243
transform 1 0 1796 0 1 675
box -3 -3 3 3
use XOR2X1  XOR2X1_34
timestamp 1524952243
transform 1 0 1760 0 -1 770
box -8 -3 64 105
use OAI21X1  OAI21X1_69
timestamp 1524952243
transform 1 0 1816 0 -1 770
box -8 -3 34 105
use AOI21X1  AOI21X1_9
timestamp 1524952243
transform 1 0 1848 0 -1 770
box -7 -3 39 105
use NOR2X1  NOR2X1_38
timestamp 1524952243
transform 1 0 1880 0 -1 770
box -8 -3 32 105
use M3_M2  M3_M2_1767
timestamp 1524952243
transform 1 0 1940 0 1 675
box -3 -3 3 3
use AOI22X1  AOI22X1_48
timestamp 1524952243
transform 1 0 1904 0 -1 770
box -8 -3 46 105
use top_module_VIA0  top_module_VIA0_25
timestamp 1524952243
transform 1 0 1994 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_1785
timestamp 1524952243
transform 1 0 172 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1524952243
transform 1 0 140 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1524952243
transform 1 0 68 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1524952243
transform 1 0 116 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1641
timestamp 1524952243
transform 1 0 68 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1524952243
transform 1 0 132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1524952243
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1524952243
transform 1 0 156 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1795
timestamp 1524952243
transform 1 0 188 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1524952243
transform 1 0 212 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_1637
timestamp 1524952243
transform 1 0 188 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_1831
timestamp 1524952243
transform 1 0 204 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1638
timestamp 1524952243
transform 1 0 220 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1524952243
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1524952243
transform 1 0 212 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1856
timestamp 1524952243
transform 1 0 220 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1646
timestamp 1524952243
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1524952243
transform 1 0 180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1524952243
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1524952243
transform 1 0 212 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1909
timestamp 1524952243
transform 1 0 212 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1524952243
transform 1 0 268 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1524952243
transform 1 0 284 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1524952243
transform 1 0 316 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1524952243
transform 1 0 260 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1647
timestamp 1524952243
transform 1 0 260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1524952243
transform 1 0 268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1524952243
transform 1 0 244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1524952243
transform 1 0 252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1524952243
transform 1 0 268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1890
timestamp 1524952243
transform 1 0 244 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1524952243
transform 1 0 268 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1524952243
transform 1 0 292 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1524952243
transform 1 0 332 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1524952243
transform 1 0 324 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1649
timestamp 1524952243
transform 1 0 292 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1857
timestamp 1524952243
transform 1 0 300 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1650
timestamp 1524952243
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1524952243
transform 1 0 324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1524952243
transform 1 0 292 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1875
timestamp 1524952243
transform 1 0 300 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1708
timestamp 1524952243
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1524952243
transform 1 0 324 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1876
timestamp 1524952243
transform 1 0 332 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1761
timestamp 1524952243
transform 1 0 284 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_1910
timestamp 1524952243
transform 1 0 276 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1524952243
transform 1 0 316 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1762
timestamp 1524952243
transform 1 0 332 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_1911
timestamp 1524952243
transform 1 0 316 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1524952243
transform 1 0 364 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1524952243
transform 1 0 452 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1524952243
transform 1 0 388 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1524952243
transform 1 0 380 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1524952243
transform 1 0 564 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1524952243
transform 1 0 476 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1524952243
transform 1 0 532 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1524952243
transform 1 0 460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1524952243
transform 1 0 588 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_1652
timestamp 1524952243
transform 1 0 388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1524952243
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1524952243
transform 1 0 460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1524952243
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1524952243
transform 1 0 348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1524952243
transform 1 0 364 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1877
timestamp 1524952243
transform 1 0 396 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1712
timestamp 1524952243
transform 1 0 452 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1893
timestamp 1524952243
transform 1 0 444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1524952243
transform 1 0 524 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1524952243
transform 1 0 556 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1524952243
transform 1 0 756 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1524952243
transform 1 0 772 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1524952243
transform 1 0 612 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1524952243
transform 1 0 644 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1524952243
transform 1 0 732 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1524952243
transform 1 0 620 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1524952243
transform 1 0 604 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1656
timestamp 1524952243
transform 1 0 564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1524952243
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1524952243
transform 1 0 588 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1861
timestamp 1524952243
transform 1 0 596 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1524952243
transform 1 0 652 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1659
timestamp 1524952243
transform 1 0 612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1524952243
transform 1 0 628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1524952243
transform 1 0 476 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1524952243
transform 1 0 564 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1894
timestamp 1524952243
transform 1 0 516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1524952243
transform 1 0 468 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1524952243
transform 1 0 572 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1524952243
transform 1 0 636 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1524952243
transform 1 0 772 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1524952243
transform 1 0 756 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1661
timestamp 1524952243
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1524952243
transform 1 0 732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1524952243
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1524952243
transform 1 0 580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1524952243
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1524952243
transform 1 0 604 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1895
timestamp 1524952243
transform 1 0 580 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1524952243
transform 1 0 564 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1524952243
transform 1 0 580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1524952243
transform 1 0 612 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1718
timestamp 1524952243
transform 1 0 620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1880
timestamp 1524952243
transform 1 0 628 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1524952243
transform 1 0 772 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1719
timestamp 1524952243
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1524952243
transform 1 0 652 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1896
timestamp 1524952243
transform 1 0 620 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1524952243
transform 1 0 732 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1721
timestamp 1524952243
transform 1 0 740 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1897
timestamp 1524952243
transform 1 0 676 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1524952243
transform 1 0 644 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1524952243
transform 1 0 876 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1524952243
transform 1 0 900 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1524952243
transform 1 0 940 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1524952243
transform 1 0 1028 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1524952243
transform 1 0 1076 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1524952243
transform 1 0 1068 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1524952243
transform 1 0 1084 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1524952243
transform 1 0 972 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1524952243
transform 1 0 988 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1524952243
transform 1 0 1028 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1524952243
transform 1 0 884 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1524952243
transform 1 0 900 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1524952243
transform 1 0 932 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1524952243
transform 1 0 1004 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1524952243
transform 1 0 844 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1524952243
transform 1 0 892 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1664
timestamp 1524952243
transform 1 0 844 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1864
timestamp 1524952243
transform 1 0 876 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1665
timestamp 1524952243
transform 1 0 884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1524952243
transform 1 0 900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1524952243
transform 1 0 916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1524952243
transform 1 0 788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1524952243
transform 1 0 804 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1524952243
transform 1 0 756 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1524952243
transform 1 0 844 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1524952243
transform 1 0 980 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1524952243
transform 1 0 1060 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1668
timestamp 1524952243
transform 1 0 964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1524952243
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1524952243
transform 1 0 1028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1524952243
transform 1 0 892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1524952243
transform 1 0 908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1524952243
transform 1 0 924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1524952243
transform 1 0 940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1898
timestamp 1524952243
transform 1 0 908 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1524952243
transform 1 0 1020 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1728
timestamp 1524952243
transform 1 0 1028 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1899
timestamp 1524952243
transform 1 0 964 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1524952243
transform 1 0 988 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1524952243
transform 1 0 956 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1524952243
transform 1 0 1140 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1524952243
transform 1 0 1204 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1524952243
transform 1 0 1188 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1524952243
transform 1 0 1156 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1524952243
transform 1 0 1132 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1524952243
transform 1 0 1100 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1524952243
transform 1 0 1140 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1524952243
transform 1 0 1100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1524952243
transform 1 0 1076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1524952243
transform 1 0 1084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1524952243
transform 1 0 1196 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1524952243
transform 1 0 1156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1524952243
transform 1 0 1188 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1823
timestamp 1524952243
transform 1 0 1220 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1674
timestamp 1524952243
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1524952243
transform 1 0 1228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1524952243
transform 1 0 1132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1524952243
transform 1 0 1140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1524952243
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1884
timestamp 1524952243
transform 1 0 1196 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1734
timestamp 1524952243
transform 1 0 1220 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1918
timestamp 1524952243
transform 1 0 1132 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1524952243
transform 1 0 1148 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1524952243
transform 1 0 1188 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1524952243
transform 1 0 1204 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1524952243
transform 1 0 1268 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_1636
timestamp 1524952243
transform 1 0 1268 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_1824
timestamp 1524952243
transform 1 0 1276 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1524952243
transform 1 0 1340 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1524952243
transform 1 0 1316 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1640
timestamp 1524952243
transform 1 0 1276 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_1844
timestamp 1524952243
transform 1 0 1284 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1524952243
transform 1 0 1292 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1524952243
transform 1 0 1348 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1676
timestamp 1524952243
transform 1 0 1316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1524952243
transform 1 0 1324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1524952243
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1885
timestamp 1524952243
transform 1 0 1268 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1736
timestamp 1524952243
transform 1 0 1276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1524952243
transform 1 0 1292 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1866
timestamp 1524952243
transform 1 0 1356 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1678
timestamp 1524952243
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1524952243
transform 1 0 1380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1524952243
transform 1 0 1356 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1886
timestamp 1524952243
transform 1 0 1364 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1739
timestamp 1524952243
transform 1 0 1380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1524952243
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1901
timestamp 1524952243
transform 1 0 1340 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1524952243
transform 1 0 1356 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1524952243
transform 1 0 1316 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1524952243
transform 1 0 1444 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1524952243
transform 1 0 1404 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1524952243
transform 1 0 1428 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1680
timestamp 1524952243
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1867
timestamp 1524952243
transform 1 0 1404 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1524952243
transform 1 0 1484 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1524952243
transform 1 0 1468 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1524952243
transform 1 0 1516 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1524952243
transform 1 0 1508 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1681
timestamp 1524952243
transform 1 0 1428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1524952243
transform 1 0 1452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1524952243
transform 1 0 1476 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1868
timestamp 1524952243
transform 1 0 1500 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1524952243
transform 1 0 1548 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1524952243
transform 1 0 1580 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1524952243
transform 1 0 1652 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1524952243
transform 1 0 1556 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1524952243
transform 1 0 1604 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1684
timestamp 1524952243
transform 1 0 1508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1524952243
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1524952243
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1524952243
transform 1 0 1404 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1887
timestamp 1524952243
transform 1 0 1452 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1742
timestamp 1524952243
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1888
timestamp 1524952243
transform 1 0 1476 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1743
timestamp 1524952243
transform 1 0 1484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1524952243
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1524952243
transform 1 0 1500 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1923
timestamp 1524952243
transform 1 0 1404 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1524952243
transform 1 0 1460 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1524952243
transform 1 0 1540 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1687
timestamp 1524952243
transform 1 0 1556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1524952243
transform 1 0 1580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1524952243
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1524952243
transform 1 0 1540 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1903
timestamp 1524952243
transform 1 0 1500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1524952243
transform 1 0 1524 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1524952243
transform 1 0 1492 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1524952243
transform 1 0 1540 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1524952243
transform 1 0 1588 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1689
timestamp 1524952243
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1524952243
transform 1 0 1604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1524952243
transform 1 0 1612 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1851
timestamp 1524952243
transform 1 0 1660 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1524952243
transform 1 0 1732 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1524952243
transform 1 0 1812 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1524952243
transform 1 0 1844 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1524952243
transform 1 0 1764 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1524952243
transform 1 0 1780 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_1690
timestamp 1524952243
transform 1 0 1668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1524952243
transform 1 0 1684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1524952243
transform 1 0 1700 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1871
timestamp 1524952243
transform 1 0 1732 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1524952243
transform 1 0 1756 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1750
timestamp 1524952243
transform 1 0 1660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1524952243
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1524952243
transform 1 0 1692 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1889
timestamp 1524952243
transform 1 0 1700 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_1753
timestamp 1524952243
transform 1 0 1708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1905
timestamp 1524952243
transform 1 0 1692 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1524952243
transform 1 0 1668 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_1754
timestamp 1524952243
transform 1 0 1756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1524952243
transform 1 0 1764 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1906
timestamp 1524952243
transform 1 0 1764 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1524952243
transform 1 0 1820 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1524952243
transform 1 0 1868 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1693
timestamp 1524952243
transform 1 0 1820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1524952243
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1524952243
transform 1 0 1836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1524952243
transform 1 0 1852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1524952243
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1524952243
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1928
timestamp 1524952243
transform 1 0 1772 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1524952243
transform 1 0 1860 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1697
timestamp 1524952243
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1524952243
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1524952243
transform 1 0 1860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1907
timestamp 1524952243
transform 1 0 1836 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1524952243
transform 1 0 1844 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1524952243
transform 1 0 1932 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1524952243
transform 1 0 1932 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1524952243
transform 1 0 1884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1524952243
transform 1 0 1916 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1698
timestamp 1524952243
transform 1 0 1908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1524952243
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_1874
timestamp 1524952243
transform 1 0 1948 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1760
timestamp 1524952243
transform 1 0 1948 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_1908
timestamp 1524952243
transform 1 0 1932 0 1 595
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_26
timestamp 1524952243
transform 1 0 48 0 1 570
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_77
timestamp 1524952243
transform -1 0 168 0 1 570
box -8 -3 104 105
use INVX2  INVX2_108
timestamp 1524952243
transform -1 0 184 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_1930
timestamp 1524952243
transform 1 0 220 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_70
timestamp 1524952243
transform -1 0 216 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1524952243
transform -1 0 248 0 1 570
box -8 -3 34 105
use INVX2  INVX2_109
timestamp 1524952243
transform 1 0 248 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_1931
timestamp 1524952243
transform 1 0 292 0 1 575
box -3 -3 3 3
use NOR2X1  NOR2X1_39
timestamp 1524952243
transform -1 0 288 0 1 570
box -8 -3 32 105
use AOI22X1  AOI22X1_49
timestamp 1524952243
transform -1 0 328 0 1 570
box -8 -3 46 105
use NOR2X1  NOR2X1_40
timestamp 1524952243
transform 1 0 328 0 1 570
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_78
timestamp 1524952243
transform 1 0 352 0 1 570
box -8 -3 104 105
use INVX2  INVX2_113
timestamp 1524952243
transform 1 0 448 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_1932
timestamp 1524952243
transform 1 0 548 0 1 575
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_81
timestamp 1524952243
transform 1 0 464 0 1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_15
timestamp 1524952243
transform 1 0 560 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1524952243
transform 1 0 600 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_1933
timestamp 1524952243
transform 1 0 652 0 1 575
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_82
timestamp 1524952243
transform 1 0 640 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_1934
timestamp 1524952243
transform 1 0 748 0 1 575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_32
timestamp 1524952243
transform -1 0 792 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_1935
timestamp 1524952243
transform 1 0 804 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1524952243
transform 1 0 884 0 1 575
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_83
timestamp 1524952243
transform 1 0 792 0 1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_17
timestamp 1524952243
transform 1 0 888 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_1937
timestamp 1524952243
transform 1 0 988 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1524952243
transform 1 0 1004 0 1 575
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_84
timestamp 1524952243
transform 1 0 928 0 1 570
box -8 -3 104 105
use XNOR2X1  XNOR2X1_33
timestamp 1524952243
transform -1 0 1080 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_1939
timestamp 1524952243
transform 1 0 1124 0 1 575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_34
timestamp 1524952243
transform -1 0 1136 0 1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_35
timestamp 1524952243
transform -1 0 1192 0 1 570
box -8 -3 64 105
use OAI21X1  OAI21X1_73
timestamp 1524952243
transform -1 0 1224 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1524952243
transform 1 0 1224 0 1 570
box -8 -3 34 105
use NAND3X1  NAND3X1_24
timestamp 1524952243
transform -1 0 1288 0 1 570
box -8 -3 40 105
use XOR2X1  XOR2X1_36
timestamp 1524952243
transform 1 0 1288 0 1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_52
timestamp 1524952243
transform 1 0 1344 0 1 570
box -8 -3 46 105
use INVX2  INVX2_115
timestamp 1524952243
transform 1 0 1384 0 1 570
box -9 -3 26 105
use XOR2X1  XOR2X1_37
timestamp 1524952243
transform 1 0 1400 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_1940
timestamp 1524952243
transform 1 0 1468 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_53
timestamp 1524952243
transform -1 0 1496 0 1 570
box -8 -3 46 105
use INVX2  INVX2_116
timestamp 1524952243
transform 1 0 1496 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_54
timestamp 1524952243
transform 1 0 1512 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_1941
timestamp 1524952243
transform 1 0 1612 0 1 575
box -3 -3 3 3
use XOR2X1  XOR2X1_38
timestamp 1524952243
transform 1 0 1552 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_1942
timestamp 1524952243
transform 1 0 1660 0 1 575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_35
timestamp 1524952243
transform -1 0 1664 0 1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_55
timestamp 1524952243
transform 1 0 1664 0 1 570
box -8 -3 46 105
use XNOR2X1  XNOR2X1_36
timestamp 1524952243
transform -1 0 1760 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_1943
timestamp 1524952243
transform 1 0 1820 0 1 575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_37
timestamp 1524952243
transform 1 0 1760 0 1 570
box -8 -3 64 105
use INVX2  INVX2_117
timestamp 1524952243
transform 1 0 1816 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_1944
timestamp 1524952243
transform 1 0 1884 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_56
timestamp 1524952243
transform 1 0 1832 0 1 570
box -8 -3 46 105
use FILL  FILL_17
timestamp 1524952243
transform 1 0 1872 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_1945
timestamp 1524952243
transform 1 0 1932 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1524952243
transform 1 0 1948 0 1 575
box -3 -3 3 3
use XOR2X1  XOR2X1_39
timestamp 1524952243
transform -1 0 1936 0 1 570
box -8 -3 64 105
use FILL  FILL_18
timestamp 1524952243
transform 1 0 1936 0 1 570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_27
timestamp 1524952243
transform 1 0 1970 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_1947
timestamp 1524952243
transform 1 0 132 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1524952243
transform 1 0 140 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1524952243
transform 1 0 188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1524952243
transform 1 0 124 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1767
timestamp 1524952243
transform 1 0 156 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2012
timestamp 1524952243
transform 1 0 172 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1768
timestamp 1524952243
transform 1 0 180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1524952243
transform 1 0 196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1524952243
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1524952243
transform 1 0 76 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1524952243
transform 1 0 132 0 1 526
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1524952243
transform 1 0 172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1524952243
transform 1 0 188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1524952243
transform 1 0 204 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2041
timestamp 1524952243
transform 1 0 108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1524952243
transform 1 0 76 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1524952243
transform 1 0 236 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1524952243
transform 1 0 228 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1524952243
transform 1 0 244 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1765
timestamp 1524952243
transform 1 0 236 0 1 536
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1524952243
transform 1 0 228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1524952243
transform 1 0 236 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2042
timestamp 1524952243
transform 1 0 204 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1524952243
transform 1 0 212 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_2098
timestamp 1524952243
transform 1 0 172 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1524952243
transform 1 0 212 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1524952243
transform 1 0 228 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1524952243
transform 1 0 228 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1524952243
transform 1 0 276 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1524952243
transform 1 0 268 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1524952243
transform 1 0 308 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_1763
timestamp 1524952243
transform 1 0 300 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1524952243
transform 1 0 268 0 1 536
box -2 -2 2 2
use M3_M2  M3_M2_2013
timestamp 1524952243
transform 1 0 276 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1524952243
transform 1 0 324 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1771
timestamp 1524952243
transform 1 0 292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1524952243
transform 1 0 308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1524952243
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1524952243
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1524952243
transform 1 0 260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1524952243
transform 1 0 276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1524952243
transform 1 0 300 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2043
timestamp 1524952243
transform 1 0 252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1524952243
transform 1 0 260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1524952243
transform 1 0 292 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1524952243
transform 1 0 268 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1524952243
transform 1 0 260 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_1844
timestamp 1524952243
transform 1 0 316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1524952243
transform 1 0 324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2044
timestamp 1524952243
transform 1 0 316 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1524952243
transform 1 0 332 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1774
timestamp 1524952243
transform 1 0 340 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2025
timestamp 1524952243
transform 1 0 332 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1846
timestamp 1524952243
transform 1 0 340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_1963
timestamp 1524952243
transform 1 0 412 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1524952243
transform 1 0 452 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1524952243
transform 1 0 444 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1775
timestamp 1524952243
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1524952243
transform 1 0 452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1524952243
transform 1 0 348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1524952243
transform 1 0 388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1524952243
transform 1 0 444 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2026
timestamp 1524952243
transform 1 0 452 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1524952243
transform 1 0 348 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1524952243
transform 1 0 388 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1524952243
transform 1 0 444 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1524952243
transform 1 0 340 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1524952243
transform 1 0 452 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1524952243
transform 1 0 396 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1524952243
transform 1 0 444 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1524952243
transform 1 0 476 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1524952243
transform 1 0 468 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1777
timestamp 1524952243
transform 1 0 468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1524952243
transform 1 0 460 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2027
timestamp 1524952243
transform 1 0 468 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1524952243
transform 1 0 500 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1524952243
transform 1 0 532 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1778
timestamp 1524952243
transform 1 0 532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1524952243
transform 1 0 548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1524952243
transform 1 0 476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1524952243
transform 1 0 484 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2028
timestamp 1524952243
transform 1 0 500 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1853
timestamp 1524952243
transform 1 0 516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2048
timestamp 1524952243
transform 1 0 484 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1524952243
transform 1 0 500 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1524952243
transform 1 0 556 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1780
timestamp 1524952243
transform 1 0 564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1524952243
transform 1 0 556 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2029
timestamp 1524952243
transform 1 0 564 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1524952243
transform 1 0 628 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1524952243
transform 1 0 676 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1524952243
transform 1 0 692 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1524952243
transform 1 0 636 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1524952243
transform 1 0 652 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1781
timestamp 1524952243
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1524952243
transform 1 0 644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1524952243
transform 1 0 652 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2016
timestamp 1524952243
transform 1 0 660 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1855
timestamp 1524952243
transform 1 0 588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1524952243
transform 1 0 620 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2049
timestamp 1524952243
transform 1 0 556 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1524952243
transform 1 0 564 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1524952243
transform 1 0 628 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1857
timestamp 1524952243
transform 1 0 636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2031
timestamp 1524952243
transform 1 0 644 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1524952243
transform 1 0 724 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1524952243
transform 1 0 748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1524952243
transform 1 0 788 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1524952243
transform 1 0 724 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1784
timestamp 1524952243
transform 1 0 716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1524952243
transform 1 0 724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1524952243
transform 1 0 652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1524952243
transform 1 0 660 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2050
timestamp 1524952243
transform 1 0 620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1524952243
transform 1 0 596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1524952243
transform 1 0 676 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1524952243
transform 1 0 732 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1786
timestamp 1524952243
transform 1 0 740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1524952243
transform 1 0 756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1524952243
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1524952243
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1524952243
transform 1 0 756 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2051
timestamp 1524952243
transform 1 0 660 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1524952243
transform 1 0 684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1524952243
transform 1 0 740 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1524952243
transform 1 0 892 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1524952243
transform 1 0 844 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1788
timestamp 1524952243
transform 1 0 804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1524952243
transform 1 0 820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1524952243
transform 1 0 852 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_1953
timestamp 1524952243
transform 1 0 980 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1524952243
transform 1 0 916 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1524952243
transform 1 0 964 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1524952243
transform 1 0 908 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1791
timestamp 1524952243
transform 1 0 900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1524952243
transform 1 0 908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1524952243
transform 1 0 804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1524952243
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1524952243
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1524952243
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1524952243
transform 1 0 900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2053
timestamp 1524952243
transform 1 0 804 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1524952243
transform 1 0 908 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1524952243
transform 1 0 1028 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1524952243
transform 1 0 1020 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1524952243
transform 1 0 956 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1524952243
transform 1 0 972 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1793
timestamp 1524952243
transform 1 0 956 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2018
timestamp 1524952243
transform 1 0 980 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1524952243
transform 1 0 1076 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1524952243
transform 1 0 1092 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1794
timestamp 1524952243
transform 1 0 1028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1524952243
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1524952243
transform 1 0 940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1524952243
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1524952243
transform 1 0 972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1524952243
transform 1 0 980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1524952243
transform 1 0 1012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1524952243
transform 1 0 1028 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1524952243
transform 1 0 884 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1524952243
transform 1 0 900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1524952243
transform 1 0 828 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1524952243
transform 1 0 852 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1524952243
transform 1 0 964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1524952243
transform 1 0 980 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1524952243
transform 1 0 916 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1524952243
transform 1 0 1028 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1796
timestamp 1524952243
transform 1 0 1092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1524952243
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2019
timestamp 1524952243
transform 1 0 1116 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1524952243
transform 1 0 1172 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1524952243
transform 1 0 1188 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1798
timestamp 1524952243
transform 1 0 1132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1524952243
transform 1 0 1140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1524952243
transform 1 0 1148 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1524952243
transform 1 0 1164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1524952243
transform 1 0 1172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1524952243
transform 1 0 1084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1524952243
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1524952243
transform 1 0 1108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2034
timestamp 1524952243
transform 1 0 1116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1524952243
transform 1 0 1084 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1524952243
transform 1 0 1108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1524952243
transform 1 0 988 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1524952243
transform 1 0 1036 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1524952243
transform 1 0 1076 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1524952243
transform 1 0 972 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1524952243
transform 1 0 1100 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1524952243
transform 1 0 1180 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1877
timestamp 1524952243
transform 1 0 1156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1524952243
transform 1 0 1172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1524952243
transform 1 0 1132 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_2061
timestamp 1524952243
transform 1 0 1140 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1524952243
transform 1 0 1172 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1524952243
transform 1 0 1140 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1524952243
transform 1 0 1164 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1524952243
transform 1 0 1220 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1524952243
transform 1 0 1212 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1524952243
transform 1 0 1236 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1524952243
transform 1 0 1260 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1524952243
transform 1 0 1204 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1803
timestamp 1524952243
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2001
timestamp 1524952243
transform 1 0 1252 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1804
timestamp 1524952243
transform 1 0 1252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1524952243
transform 1 0 1260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1524952243
transform 1 0 1196 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2035
timestamp 1524952243
transform 1 0 1220 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1880
timestamp 1524952243
transform 1 0 1260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1524952243
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1524952243
transform 1 0 1292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_1981
timestamp 1524952243
transform 1 0 1324 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1524952243
transform 1 0 1372 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1524952243
transform 1 0 1364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1524952243
transform 1 0 1348 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1764
timestamp 1524952243
transform 1 0 1356 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_2003
timestamp 1524952243
transform 1 0 1380 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1806
timestamp 1524952243
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2021
timestamp 1524952243
transform 1 0 1332 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1807
timestamp 1524952243
transform 1 0 1340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1524952243
transform 1 0 1348 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2022
timestamp 1524952243
transform 1 0 1356 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1809
timestamp 1524952243
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1524952243
transform 1 0 1372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1524952243
transform 1 0 1332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1524952243
transform 1 0 1196 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_2062
timestamp 1524952243
transform 1 0 1236 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1524952243
transform 1 0 1260 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1524952243
transform 1 0 1292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1524952243
transform 1 0 1308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1524952243
transform 1 0 1220 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1524952243
transform 1 0 1284 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1524952243
transform 1 0 1316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1524952243
transform 1 0 1308 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1524952243
transform 1 0 1324 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1524952243
transform 1 0 1436 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1524952243
transform 1 0 1460 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1524952243
transform 1 0 1428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1811
timestamp 1524952243
transform 1 0 1428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1524952243
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1524952243
transform 1 0 1380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1524952243
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2036
timestamp 1524952243
transform 1 0 1404 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1813
timestamp 1524952243
transform 1 0 1484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1524952243
transform 1 0 1492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1524952243
transform 1 0 1508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1524952243
transform 1 0 1516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1524952243
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1524952243
transform 1 0 1436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1524952243
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1524952243
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2066
timestamp 1524952243
transform 1 0 1396 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1524952243
transform 1 0 1428 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1524952243
transform 1 0 1396 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1524952243
transform 1 0 1420 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1524952243
transform 1 0 1436 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_1889
timestamp 1524952243
transform 1 0 1508 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2037
timestamp 1524952243
transform 1 0 1516 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1524952243
transform 1 0 1604 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1818
timestamp 1524952243
transform 1 0 1596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1524952243
transform 1 0 1604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1524952243
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1524952243
transform 1 0 1548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1524952243
transform 1 0 1572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1524952243
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2092
timestamp 1524952243
transform 1 0 1508 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1524952243
transform 1 0 1604 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1524952243
transform 1 0 1548 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1524952243
transform 1 0 1596 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1524952243
transform 1 0 1540 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1524952243
transform 1 0 1572 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1524952243
transform 1 0 1492 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1524952243
transform 1 0 1516 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1524952243
transform 1 0 1460 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1524952243
transform 1 0 1580 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1524952243
transform 1 0 1564 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1524952243
transform 1 0 1652 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1524952243
transform 1 0 1684 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1524952243
transform 1 0 1708 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1820
timestamp 1524952243
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1524952243
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1524952243
transform 1 0 1684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1524952243
transform 1 0 1700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1524952243
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2095
timestamp 1524952243
transform 1 0 1652 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1524952243
transform 1 0 1748 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1524952243
transform 1 0 1748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1524952243
transform 1 0 1724 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2113
timestamp 1524952243
transform 1 0 1756 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1524952243
transform 1 0 1692 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1524952243
transform 1 0 1724 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1524952243
transform 1 0 1756 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1524952243
transform 1 0 1764 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1825
timestamp 1524952243
transform 1 0 1764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1524952243
transform 1 0 1772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1524952243
transform 1 0 1764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1524952243
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_1985
timestamp 1524952243
transform 1 0 1820 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1827
timestamp 1524952243
transform 1 0 1796 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2023
timestamp 1524952243
transform 1 0 1804 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1828
timestamp 1524952243
transform 1 0 1812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1524952243
transform 1 0 1820 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2024
timestamp 1524952243
transform 1 0 1828 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1898
timestamp 1524952243
transform 1 0 1780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1524952243
transform 1 0 1788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2039
timestamp 1524952243
transform 1 0 1796 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1900
timestamp 1524952243
transform 1 0 1804 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2040
timestamp 1524952243
transform 1 0 1812 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1901
timestamp 1524952243
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1524952243
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2070
timestamp 1524952243
transform 1 0 1788 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1524952243
transform 1 0 1812 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1524952243
transform 1 0 1828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1524952243
transform 1 0 1820 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1524952243
transform 1 0 1796 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1524952243
transform 1 0 1876 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1524952243
transform 1 0 1876 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1830
timestamp 1524952243
transform 1 0 1876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1524952243
transform 1 0 1884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1524952243
transform 1 0 1900 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1524952243
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_2073
timestamp 1524952243
transform 1 0 1916 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1524952243
transform 1 0 1932 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1524952243
transform 1 0 2012 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1832
timestamp 1524952243
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_2115
timestamp 1524952243
transform 1 0 2012 0 1 495
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_28
timestamp 1524952243
transform 1 0 24 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_2127
timestamp 1524952243
transform 1 0 116 0 1 475
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_79
timestamp 1524952243
transform -1 0 168 0 -1 570
box -8 -3 104 105
use AOI22X1  AOI22X1_50
timestamp 1524952243
transform -1 0 208 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_2128
timestamp 1524952243
transform 1 0 220 0 1 475
box -3 -3 3 3
use OAI21X1  OAI21X1_72
timestamp 1524952243
transform -1 0 240 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_110
timestamp 1524952243
transform 1 0 240 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_51
timestamp 1524952243
transform -1 0 296 0 -1 570
box -8 -3 46 105
use NOR2X1  NOR2X1_41
timestamp 1524952243
transform 1 0 296 0 -1 570
box -8 -3 32 105
use INVX2  INVX2_111
timestamp 1524952243
transform 1 0 320 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1524952243
transform 1 0 336 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_2129
timestamp 1524952243
transform 1 0 436 0 1 475
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_80
timestamp 1524952243
transform 1 0 352 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_114
timestamp 1524952243
transform 1 0 448 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1524952243
transform 1 0 464 0 -1 570
box -9 -3 26 105
use XNOR2X1  XNOR2X1_38
timestamp 1524952243
transform 1 0 480 0 -1 570
box -8 -3 64 105
use NOR2X1  NOR2X1_42
timestamp 1524952243
transform 1 0 536 0 -1 570
box -8 -3 32 105
use XOR2X1  XOR2X1_40
timestamp 1524952243
transform 1 0 560 0 -1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_57
timestamp 1524952243
transform -1 0 656 0 -1 570
box -8 -3 46 105
use XNOR2X1  XNOR2X1_39
timestamp 1524952243
transform -1 0 712 0 -1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_58
timestamp 1524952243
transform 1 0 712 0 -1 570
box -8 -3 46 105
use XOR2X1  XOR2X1_41
timestamp 1524952243
transform -1 0 808 0 -1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_59
timestamp 1524952243
transform 1 0 808 0 -1 570
box -8 -3 46 105
use XNOR2X1  XNOR2X1_40
timestamp 1524952243
transform 1 0 848 0 -1 570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_41
timestamp 1524952243
transform 1 0 904 0 -1 570
box -8 -3 64 105
use INVX2  INVX2_119
timestamp 1524952243
transform -1 0 976 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_2130
timestamp 1524952243
transform 1 0 1028 0 1 475
box -3 -3 3 3
use XNOR2X1  XNOR2X1_42
timestamp 1524952243
transform 1 0 976 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_42
timestamp 1524952243
transform -1 0 1088 0 -1 570
box -8 -3 64 105
use INVX2  INVX2_120
timestamp 1524952243
transform 1 0 1088 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_2131
timestamp 1524952243
transform 1 0 1148 0 1 475
box -3 -3 3 3
use OAI21X1  OAI21X1_75
timestamp 1524952243
transform 1 0 1104 0 -1 570
box -8 -3 34 105
use AOI22X1  AOI22X1_60
timestamp 1524952243
transform -1 0 1176 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_2132
timestamp 1524952243
transform 1 0 1188 0 1 475
box -3 -3 3 3
use NAND2X1  NAND2X1_41
timestamp 1524952243
transform 1 0 1176 0 -1 570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_43
timestamp 1524952243
transform 1 0 1200 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_43
timestamp 1524952243
transform 1 0 1256 0 -1 570
box -8 -3 64 105
use AOI22X1  AOI22X1_61
timestamp 1524952243
transform 1 0 1312 0 -1 570
box -8 -3 46 105
use NOR2X1  NOR2X1_43
timestamp 1524952243
transform 1 0 1352 0 -1 570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_44
timestamp 1524952243
transform -1 0 1432 0 -1 570
box -8 -3 64 105
use M3_M2  M3_M2_2133
timestamp 1524952243
transform 1 0 1468 0 1 475
box -3 -3 3 3
use XOR2X1  XOR2X1_44
timestamp 1524952243
transform 1 0 1432 0 -1 570
box -8 -3 64 105
use INVX2  INVX2_121
timestamp 1524952243
transform 1 0 1488 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_2134
timestamp 1524952243
transform 1 0 1524 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_62
timestamp 1524952243
transform 1 0 1504 0 -1 570
box -8 -3 46 105
use XOR2X1  XOR2X1_45
timestamp 1524952243
transform 1 0 1544 0 -1 570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_45
timestamp 1524952243
transform -1 0 1656 0 -1 570
box -8 -3 64 105
use M3_M2  M3_M2_2135
timestamp 1524952243
transform 1 0 1684 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_63
timestamp 1524952243
transform 1 0 1656 0 -1 570
box -8 -3 46 105
use XOR2X1  XOR2X1_46
timestamp 1524952243
transform -1 0 1752 0 -1 570
box -8 -3 64 105
use M3_M2  M3_M2_2136
timestamp 1524952243
transform 1 0 1772 0 1 475
box -3 -3 3 3
use INVX2  INVX2_122
timestamp 1524952243
transform -1 0 1768 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1524952243
transform 1 0 1768 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_2137
timestamp 1524952243
transform 1 0 1828 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_64
timestamp 1524952243
transform -1 0 1824 0 -1 570
box -8 -3 46 105
use XNOR2X1  XNOR2X1_46
timestamp 1524952243
transform -1 0 1880 0 -1 570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_47
timestamp 1524952243
transform -1 0 1936 0 -1 570
box -8 -3 64 105
use FILL  FILL_19
timestamp 1524952243
transform 1 0 1936 0 -1 570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_29
timestamp 1524952243
transform 1 0 1994 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_2138
timestamp 1524952243
transform 1 0 84 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1524952243
transform 1 0 156 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1524952243
transform 1 0 156 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1920
timestamp 1524952243
transform 1 0 76 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1524952243
transform 1 0 124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1524952243
transform 1 0 156 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2295
timestamp 1524952243
transform 1 0 76 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1524952243
transform 1 0 196 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1524952243
transform 1 0 196 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1524952243
transform 1 0 180 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1524952243
transform 1 0 292 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1524952243
transform 1 0 332 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1524952243
transform 1 0 324 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1524952243
transform 1 0 380 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1524952243
transform 1 0 468 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1524952243
transform 1 0 444 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1524952243
transform 1 0 476 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1524952243
transform 1 0 412 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1524952243
transform 1 0 316 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1524952243
transform 1 0 356 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1524952243
transform 1 0 404 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1524952243
transform 1 0 476 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1524952243
transform 1 0 444 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1524952243
transform 1 0 532 0 1 455
box -2 -2 2 2
use M3_M2  M3_M2_2162
timestamp 1524952243
transform 1 0 524 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_1910
timestamp 1524952243
transform 1 0 532 0 1 445
box -2 -2 2 2
use M3_M2  M3_M2_2182
timestamp 1524952243
transform 1 0 508 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1913
timestamp 1524952243
transform 1 0 476 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1524952243
transform 1 0 204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1524952243
transform 1 0 260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1524952243
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1524952243
transform 1 0 284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1524952243
transform 1 0 300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1524952243
transform 1 0 316 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2232
timestamp 1524952243
transform 1 0 332 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1928
timestamp 1524952243
transform 1 0 356 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2233
timestamp 1524952243
transform 1 0 364 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1929
timestamp 1524952243
transform 1 0 412 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1524952243
transform 1 0 420 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1930
timestamp 1524952243
transform 1 0 444 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2235
timestamp 1524952243
transform 1 0 452 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1524952243
transform 1 0 492 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1914
timestamp 1524952243
transform 1 0 500 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1524952243
transform 1 0 468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1524952243
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1524952243
transform 1 0 492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1524952243
transform 1 0 180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1524952243
transform 1 0 268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1524952243
transform 1 0 292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1524952243
transform 1 0 300 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2270
timestamp 1524952243
transform 1 0 180 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1524952243
transform 1 0 196 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1524952243
transform 1 0 260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1524952243
transform 1 0 212 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1524952243
transform 1 0 308 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1996
timestamp 1524952243
transform 1 0 332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2254
timestamp 1524952243
transform 1 0 356 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1524952243
transform 1 0 380 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1524952243
transform 1 0 412 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1997
timestamp 1524952243
transform 1 0 420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2274
timestamp 1524952243
transform 1 0 420 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1524952243
transform 1 0 332 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1524952243
transform 1 0 396 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1524952243
transform 1 0 468 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1524952243
transform 1 0 524 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1934
timestamp 1524952243
transform 1 0 516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1524952243
transform 1 0 500 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2275
timestamp 1524952243
transform 1 0 500 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1524952243
transform 1 0 532 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1999
timestamp 1524952243
transform 1 0 524 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1524952243
transform 1 0 532 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2299
timestamp 1524952243
transform 1 0 508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1524952243
transform 1 0 548 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1524952243
transform 1 0 548 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1524952243
transform 1 0 564 0 1 465
box -3 -3 3 3
use M2_M1  M2_M1_1909
timestamp 1524952243
transform 1 0 556 0 1 455
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1524952243
transform 1 0 556 0 1 445
box -2 -2 2 2
use M3_M2  M3_M2_2183
timestamp 1524952243
transform 1 0 556 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1524952243
transform 1 0 548 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1524952243
transform 1 0 588 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1524952243
transform 1 0 564 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1524952243
transform 1 0 644 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1524952243
transform 1 0 612 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1524952243
transform 1 0 604 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1935
timestamp 1524952243
transform 1 0 564 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2237
timestamp 1524952243
transform 1 0 572 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1936
timestamp 1524952243
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1524952243
transform 1 0 596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1524952243
transform 1 0 604 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2258
timestamp 1524952243
transform 1 0 564 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_2001
timestamp 1524952243
transform 1 0 572 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2259
timestamp 1524952243
transform 1 0 580 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_2002
timestamp 1524952243
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1524952243
transform 1 0 596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2277
timestamp 1524952243
transform 1 0 596 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1524952243
transform 1 0 676 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1524952243
transform 1 0 716 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1524952243
transform 1 0 788 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1524952243
transform 1 0 748 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1524952243
transform 1 0 708 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1524952243
transform 1 0 724 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1939
timestamp 1524952243
transform 1 0 660 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2238
timestamp 1524952243
transform 1 0 684 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1940
timestamp 1524952243
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1524952243
transform 1 0 716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1524952243
transform 1 0 652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1524952243
transform 1 0 660 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2239
timestamp 1524952243
transform 1 0 724 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1942
timestamp 1524952243
transform 1 0 732 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2240
timestamp 1524952243
transform 1 0 740 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1524952243
transform 1 0 812 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1524952243
transform 1 0 772 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1524952243
transform 1 0 804 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1943
timestamp 1524952243
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1524952243
transform 1 0 772 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1524952243
transform 1 0 788 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1524952243
transform 1 0 908 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1524952243
transform 1 0 852 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1524952243
transform 1 0 884 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1524952243
transform 1 0 916 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1524952243
transform 1 0 964 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1945
timestamp 1524952243
transform 1 0 804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1524952243
transform 1 0 812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1524952243
transform 1 0 828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1524952243
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1524952243
transform 1 0 876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1524952243
transform 1 0 884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1524952243
transform 1 0 724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1524952243
transform 1 0 740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2278
timestamp 1524952243
transform 1 0 660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1524952243
transform 1 0 708 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1524952243
transform 1 0 756 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1524952243
transform 1 0 748 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1524952243
transform 1 0 644 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1524952243
transform 1 0 660 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1524952243
transform 1 0 692 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1524952243
transform 1 0 716 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1524952243
transform 1 0 740 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_2008
timestamp 1524952243
transform 1 0 820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1524952243
transform 1 0 852 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2305
timestamp 1524952243
transform 1 0 820 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1524952243
transform 1 0 900 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1524952243
transform 1 0 940 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1524952243
transform 1 0 956 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1524952243
transform 1 0 996 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1524952243
transform 1 0 1028 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1524952243
transform 1 0 1020 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1951
timestamp 1524952243
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1524952243
transform 1 0 980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1524952243
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1524952243
transform 1 0 1012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1524952243
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1524952243
transform 1 0 908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1524952243
transform 1 0 956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1524952243
transform 1 0 972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1524952243
transform 1 0 980 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2261
timestamp 1524952243
transform 1 0 996 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_2014
timestamp 1524952243
transform 1 0 1004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1524952243
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2281
timestamp 1524952243
transform 1 0 972 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1524952243
transform 1 0 1004 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1524952243
transform 1 0 956 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_2016
timestamp 1524952243
transform 1 0 1036 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2147
timestamp 1524952243
transform 1 0 1060 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1524952243
transform 1 0 1140 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1524952243
transform 1 0 1156 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1524952243
transform 1 0 1092 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1524952243
transform 1 0 1108 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1524952243
transform 1 0 1100 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1524952243
transform 1 0 1116 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1524952243
transform 1 0 1084 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1915
timestamp 1524952243
transform 1 0 1100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1524952243
transform 1 0 1052 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1524952243
transform 1 0 1076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1524952243
transform 1 0 1084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1524952243
transform 1 0 1052 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1524952243
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1524952243
transform 1 0 1076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1524952243
transform 1 0 1052 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_2283
timestamp 1524952243
transform 1 0 1068 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1524952243
transform 1 0 1076 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1524952243
transform 1 0 1100 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1524952243
transform 1 0 1180 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1524952243
transform 1 0 1196 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1524952243
transform 1 0 1156 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1524952243
transform 1 0 1172 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_1916
timestamp 1524952243
transform 1 0 1132 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_2218
timestamp 1524952243
transform 1 0 1140 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1524952243
transform 1 0 1156 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1959
timestamp 1524952243
transform 1 0 1116 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2246
timestamp 1524952243
transform 1 0 1132 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1524952243
transform 1 0 1212 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1524952243
transform 1 0 1228 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_1960
timestamp 1524952243
transform 1 0 1140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1524952243
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1524952243
transform 1 0 1188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1524952243
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1524952243
transform 1 0 1212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1524952243
transform 1 0 1100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1524952243
transform 1 0 1108 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2262
timestamp 1524952243
transform 1 0 1116 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1524952243
transform 1 0 1100 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1524952243
transform 1 0 1220 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1524952243
transform 1 0 1308 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1524952243
transform 1 0 1324 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1524952243
transform 1 0 1252 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1524952243
transform 1 0 1268 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1524952243
transform 1 0 1284 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1965
timestamp 1524952243
transform 1 0 1236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1524952243
transform 1 0 1260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1524952243
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2263
timestamp 1524952243
transform 1 0 1188 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_2022
timestamp 1524952243
transform 1 0 1196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1524952243
transform 1 0 1220 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1524952243
transform 1 0 1228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2264
timestamp 1524952243
transform 1 0 1236 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1912
timestamp 1524952243
transform 1 0 1324 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1524952243
transform 1 0 1316 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_2248
timestamp 1524952243
transform 1 0 1300 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1968
timestamp 1524952243
transform 1 0 1308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1524952243
transform 1 0 1284 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2285
timestamp 1524952243
transform 1 0 1196 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1524952243
transform 1 0 1220 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1524952243
transform 1 0 1284 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1524952243
transform 1 0 1348 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1524952243
transform 1 0 1412 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1524952243
transform 1 0 1404 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1524952243
transform 1 0 1420 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1918
timestamp 1524952243
transform 1 0 1348 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_2223
timestamp 1524952243
transform 1 0 1372 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1524952243
transform 1 0 1388 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1524952243
transform 1 0 1404 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1919
timestamp 1524952243
transform 1 0 1412 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1524952243
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1524952243
transform 1 0 1372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1524952243
transform 1 0 1316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1524952243
transform 1 0 1332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2194
timestamp 1524952243
transform 1 0 1468 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1524952243
transform 1 0 1436 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1524952243
transform 1 0 1508 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1524952243
transform 1 0 1532 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1971
timestamp 1524952243
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1524952243
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1524952243
transform 1 0 1460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1524952243
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1524952243
transform 1 0 1484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1524952243
transform 1 0 1500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1524952243
transform 1 0 1516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1524952243
transform 1 0 1524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1524952243
transform 1 0 1556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1524952243
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1524952243
transform 1 0 1580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1524952243
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1524952243
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2265
timestamp 1524952243
transform 1 0 1460 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1524952243
transform 1 0 1436 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_2030
timestamp 1524952243
transform 1 0 1492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1524952243
transform 1 0 1508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1524952243
transform 1 0 1516 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2289
timestamp 1524952243
transform 1 0 1484 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1524952243
transform 1 0 1604 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1524952243
transform 1 0 1676 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1524952243
transform 1 0 1708 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1524952243
transform 1 0 1700 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1524952243
transform 1 0 1692 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1982
timestamp 1524952243
transform 1 0 1604 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2249
timestamp 1524952243
transform 1 0 1652 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1524952243
transform 1 0 1668 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1983
timestamp 1524952243
transform 1 0 1676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1524952243
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1524952243
transform 1 0 1588 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2266
timestamp 1524952243
transform 1 0 1596 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1524952243
transform 1 0 1588 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1524952243
transform 1 0 1580 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_2034
timestamp 1524952243
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1524952243
transform 1 0 1660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1524952243
transform 1 0 1668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1524952243
transform 1 0 1684 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2291
timestamp 1524952243
transform 1 0 1668 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1524952243
transform 1 0 1780 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1524952243
transform 1 0 1764 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1524952243
transform 1 0 1748 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1524952243
transform 1 0 1764 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1524952243
transform 1 0 1788 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1524952243
transform 1 0 1732 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1524952243
transform 1 0 1780 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1985
timestamp 1524952243
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1524952243
transform 1 0 1756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1524952243
transform 1 0 1764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1524952243
transform 1 0 1708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2252
timestamp 1524952243
transform 1 0 1796 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_2039
timestamp 1524952243
transform 1 0 1756 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2267
timestamp 1524952243
transform 1 0 1764 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1524952243
transform 1 0 1716 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1988
timestamp 1524952243
transform 1 0 1836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1524952243
transform 1 0 1812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1524952243
transform 1 0 1820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1524952243
transform 1 0 1828 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2268
timestamp 1524952243
transform 1 0 1836 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1524952243
transform 1 0 1884 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1524952243
transform 1 0 1916 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_1989
timestamp 1524952243
transform 1 0 1884 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2253
timestamp 1524952243
transform 1 0 1892 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_2043
timestamp 1524952243
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1524952243
transform 1 0 1852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1524952243
transform 1 0 1860 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_2292
timestamp 1524952243
transform 1 0 1812 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1524952243
transform 1 0 1844 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1524952243
transform 1 0 1780 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1524952243
transform 1 0 1916 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_2047
timestamp 1524952243
transform 1 0 1916 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_2311
timestamp 1524952243
transform 1 0 1852 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1524952243
transform 1 0 1892 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1990
timestamp 1524952243
transform 1 0 1932 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_2294
timestamp 1524952243
transform 1 0 1940 0 1 395
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_30
timestamp 1524952243
transform 1 0 48 0 1 370
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_85
timestamp 1524952243
transform -1 0 168 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_2313
timestamp 1524952243
transform 1 0 244 0 1 375
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_86
timestamp 1524952243
transform 1 0 168 0 1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_65
timestamp 1524952243
transform -1 0 304 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_2314
timestamp 1524952243
transform 1 0 324 0 1 375
box -3 -3 3 3
use INVX2  INVX2_124
timestamp 1524952243
transform 1 0 304 0 1 370
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_87
timestamp 1524952243
transform 1 0 320 0 1 370
box -8 -3 104 105
use XOR2X1  XOR2X1_47
timestamp 1524952243
transform 1 0 416 0 1 370
box -8 -3 64 105
use NAND2X1  NAND2X1_42
timestamp 1524952243
transform -1 0 496 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_76
timestamp 1524952243
transform -1 0 528 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_2315
timestamp 1524952243
transform 1 0 540 0 1 375
box -3 -3 3 3
use FILL  FILL_20
timestamp 1524952243
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_21
timestamp 1524952243
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_22
timestamp 1524952243
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_23
timestamp 1524952243
transform 1 0 552 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_66
timestamp 1524952243
transform -1 0 600 0 1 370
box -8 -3 46 105
use XNOR2X1  XNOR2X1_48
timestamp 1524952243
transform -1 0 656 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_48
timestamp 1524952243
transform -1 0 712 0 1 370
box -8 -3 64 105
use AOI22X1  AOI22X1_67
timestamp 1524952243
transform -1 0 752 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_2316
timestamp 1524952243
transform 1 0 780 0 1 375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_49
timestamp 1524952243
transform -1 0 808 0 1 370
box -8 -3 64 105
use AOI22X1  AOI22X1_68
timestamp 1524952243
transform 1 0 808 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_2317
timestamp 1524952243
transform 1 0 860 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_49
timestamp 1524952243
transform 1 0 848 0 1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_50
timestamp 1524952243
transform -1 0 960 0 1 370
box -8 -3 64 105
use INVX2  INVX2_125
timestamp 1524952243
transform -1 0 976 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_2318
timestamp 1524952243
transform 1 0 996 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_69
timestamp 1524952243
transform 1 0 976 0 1 370
box -8 -3 46 105
use FILL  FILL_24
timestamp 1524952243
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_25
timestamp 1524952243
transform 1 0 1024 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_2319
timestamp 1524952243
transform 1 0 1060 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1524952243
transform 1 0 1076 0 1 375
box -3 -3 3 3
use NOR2X1  NOR2X1_44
timestamp 1524952243
transform -1 0 1056 0 1 370
box -8 -3 32 105
use INVX2  INVX2_126
timestamp 1524952243
transform -1 0 1072 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_2321
timestamp 1524952243
transform 1 0 1108 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_77
timestamp 1524952243
transform 1 0 1072 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1524952243
transform 1 0 1104 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_2322
timestamp 1524952243
transform 1 0 1164 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1524952243
transform 1 0 1180 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_50
timestamp 1524952243
transform 1 0 1136 0 1 370
box -8 -3 64 105
use M3_M2  M3_M2_2324
timestamp 1524952243
transform 1 0 1204 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_70
timestamp 1524952243
transform 1 0 1192 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_2325
timestamp 1524952243
transform 1 0 1268 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_51
timestamp 1524952243
transform 1 0 1232 0 1 370
box -8 -3 64 105
use AND2X2  AND2X2_22
timestamp 1524952243
transform -1 0 1320 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1524952243
transform 1 0 1320 0 1 370
box -8 -3 40 105
use XOR2X1  XOR2X1_52
timestamp 1524952243
transform -1 0 1408 0 1 370
box -8 -3 64 105
use OAI21X1  OAI21X1_79
timestamp 1524952243
transform -1 0 1440 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_2326
timestamp 1524952243
transform 1 0 1468 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_71
timestamp 1524952243
transform 1 0 1440 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1524952243
transform 1 0 1480 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_2327
timestamp 1524952243
transform 1 0 1532 0 1 375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_51
timestamp 1524952243
transform 1 0 1520 0 1 370
box -8 -3 64 105
use FILL  FILL_26
timestamp 1524952243
transform 1 0 1576 0 1 370
box -8 -3 16 105
use INVX2  INVX2_127
timestamp 1524952243
transform 1 0 1584 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_2328
timestamp 1524952243
transform 1 0 1636 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1524952243
transform 1 0 1660 0 1 375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_52
timestamp 1524952243
transform 1 0 1600 0 1 370
box -8 -3 64 105
use AOI22X1  AOI22X1_73
timestamp 1524952243
transform -1 0 1696 0 1 370
box -8 -3 46 105
use FILL  FILL_27
timestamp 1524952243
transform 1 0 1696 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_2330
timestamp 1524952243
transform 1 0 1764 0 1 375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_53
timestamp 1524952243
transform 1 0 1704 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_53
timestamp 1524952243
transform 1 0 1760 0 1 370
box -8 -3 64 105
use AOI22X1  AOI22X1_74
timestamp 1524952243
transform 1 0 1816 0 1 370
box -8 -3 46 105
use XOR2X1  XOR2X1_54
timestamp 1524952243
transform 1 0 1856 0 1 370
box -8 -3 64 105
use NOR2X1  NOR2X1_45
timestamp 1524952243
transform 1 0 1912 0 1 370
box -8 -3 32 105
use FILL  FILL_28
timestamp 1524952243
transform 1 0 1936 0 1 370
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_31
timestamp 1524952243
transform 1 0 1970 0 1 370
box -10 -3 10 3
use M3_M2  M3_M2_2331
timestamp 1524952243
transform 1 0 68 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_2107
timestamp 1524952243
transform 1 0 68 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2353
timestamp 1524952243
transform 1 0 140 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1524952243
transform 1 0 148 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2053
timestamp 1524952243
transform 1 0 172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1524952243
transform 1 0 148 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2332
timestamp 1524952243
transform 1 0 268 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1524952243
transform 1 0 252 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1524952243
transform 1 0 308 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1524952243
transform 1 0 268 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1524952243
transform 1 0 292 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2054
timestamp 1524952243
transform 1 0 204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1524952243
transform 1 0 228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1524952243
transform 1 0 236 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1524952243
transform 1 0 260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1524952243
transform 1 0 268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1524952243
transform 1 0 292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1524952243
transform 1 0 300 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2406
timestamp 1524952243
transform 1 0 204 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2109
timestamp 1524952243
transform 1 0 220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1524952243
transform 1 0 204 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2407
timestamp 1524952243
transform 1 0 236 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2110
timestamp 1524952243
transform 1 0 252 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2408
timestamp 1524952243
transform 1 0 268 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2111
timestamp 1524952243
transform 1 0 292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1524952243
transform 1 0 236 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2445
timestamp 1524952243
transform 1 0 220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1524952243
transform 1 0 252 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_2162
timestamp 1524952243
transform 1 0 268 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2409
timestamp 1524952243
transform 1 0 300 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2048
timestamp 1524952243
transform 1 0 332 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1524952243
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1524952243
transform 1 0 300 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2427
timestamp 1524952243
transform 1 0 316 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1524952243
transform 1 0 292 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1524952243
transform 1 0 260 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1524952243
transform 1 0 332 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1524952243
transform 1 0 332 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1524952243
transform 1 0 404 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1524952243
transform 1 0 428 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1524952243
transform 1 0 348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1524952243
transform 1 0 372 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2061
timestamp 1524952243
transform 1 0 348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1524952243
transform 1 0 372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1524952243
transform 1 0 348 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2428
timestamp 1524952243
transform 1 0 356 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1524952243
transform 1 0 420 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1524952243
transform 1 0 460 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1524952243
transform 1 0 492 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1524952243
transform 1 0 484 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2063
timestamp 1524952243
transform 1 0 420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1524952243
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1524952243
transform 1 0 460 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2397
timestamp 1524952243
transform 1 0 468 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2066
timestamp 1524952243
transform 1 0 484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1524952243
transform 1 0 388 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2410
timestamp 1524952243
transform 1 0 404 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2115
timestamp 1524952243
transform 1 0 420 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2411
timestamp 1524952243
transform 1 0 428 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2116
timestamp 1524952243
transform 1 0 444 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2412
timestamp 1524952243
transform 1 0 452 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2117
timestamp 1524952243
transform 1 0 476 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1524952243
transform 1 0 372 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1524952243
transform 1 0 420 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1524952243
transform 1 0 388 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_2164
timestamp 1524952243
transform 1 0 460 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2449
timestamp 1524952243
transform 1 0 460 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1524952243
transform 1 0 444 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1524952243
transform 1 0 460 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1524952243
transform 1 0 492 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2118
timestamp 1524952243
transform 1 0 500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1524952243
transform 1 0 492 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2382
timestamp 1524952243
transform 1 0 524 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2166
timestamp 1524952243
transform 1 0 516 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1524952243
transform 1 0 492 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_2450
timestamp 1524952243
transform 1 0 500 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1524952243
transform 1 0 516 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1524952243
transform 1 0 492 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1524952243
transform 1 0 556 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1524952243
transform 1 0 588 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1524952243
transform 1 0 564 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2067
timestamp 1524952243
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1524952243
transform 1 0 532 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2469
timestamp 1524952243
transform 1 0 532 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_2068
timestamp 1524952243
transform 1 0 580 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2339
timestamp 1524952243
transform 1 0 652 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1524952243
transform 1 0 700 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1524952243
transform 1 0 636 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2069
timestamp 1524952243
transform 1 0 636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1524952243
transform 1 0 700 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1524952243
transform 1 0 588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2414
timestamp 1524952243
transform 1 0 604 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2121
timestamp 1524952243
transform 1 0 620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1524952243
transform 1 0 636 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1524952243
transform 1 0 644 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1524952243
transform 1 0 668 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1524952243
transform 1 0 676 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2429
timestamp 1524952243
transform 1 0 588 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1524952243
transform 1 0 588 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1524952243
transform 1 0 732 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1524952243
transform 1 0 756 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1524952243
transform 1 0 716 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2070
timestamp 1524952243
transform 1 0 716 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2417
timestamp 1524952243
transform 1 0 708 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2124
timestamp 1524952243
transform 1 0 716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1524952243
transform 1 0 724 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2430
timestamp 1524952243
transform 1 0 700 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1524952243
transform 1 0 772 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2071
timestamp 1524952243
transform 1 0 772 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2343
timestamp 1524952243
transform 1 0 796 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1524952243
transform 1 0 788 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1524952243
transform 1 0 836 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1524952243
transform 1 0 860 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1524952243
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1524952243
transform 1 0 828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1524952243
transform 1 0 788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2431
timestamp 1524952243
transform 1 0 780 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1524952243
transform 1 0 796 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2127
timestamp 1524952243
transform 1 0 812 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2419
timestamp 1524952243
transform 1 0 820 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2128
timestamp 1524952243
transform 1 0 828 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1524952243
transform 1 0 844 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2452
timestamp 1524952243
transform 1 0 788 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1524952243
transform 1 0 828 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1524952243
transform 1 0 820 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1524952243
transform 1 0 828 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1524952243
transform 1 0 844 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1524952243
transform 1 0 860 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1524952243
transform 1 0 884 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1524952243
transform 1 0 876 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1524952243
transform 1 0 980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1524952243
transform 1 0 1004 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2074
timestamp 1524952243
transform 1 0 956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1524952243
transform 1 0 964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1524952243
transform 1 0 900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1524952243
transform 1 0 908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1524952243
transform 1 0 932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1524952243
transform 1 0 940 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2472
timestamp 1524952243
transform 1 0 892 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1524952243
transform 1 0 908 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1524952243
transform 1 0 924 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1524952243
transform 1 0 940 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1524952243
transform 1 0 932 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1524952243
transform 1 0 948 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1524952243
transform 1 0 940 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1524952243
transform 1 0 916 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1524952243
transform 1 0 1036 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1524952243
transform 1 0 1028 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2076
timestamp 1524952243
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2420
timestamp 1524952243
transform 1 0 980 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1524952243
transform 1 0 1124 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1524952243
transform 1 0 1092 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2077
timestamp 1524952243
transform 1 0 1068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1524952243
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1524952243
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1524952243
transform 1 0 1044 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2457
timestamp 1524952243
transform 1 0 980 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1524952243
transform 1 0 1052 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1524952243
transform 1 0 1044 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1524952243
transform 1 0 1124 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2079
timestamp 1524952243
transform 1 0 1124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1524952243
transform 1 0 1108 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2361
timestamp 1524952243
transform 1 0 1140 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2137
timestamp 1524952243
transform 1 0 1132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2362
timestamp 1524952243
transform 1 0 1156 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1524952243
transform 1 0 1156 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2080
timestamp 1524952243
transform 1 0 1148 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2458
timestamp 1524952243
transform 1 0 1140 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_2167
timestamp 1524952243
transform 1 0 1164 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2363
timestamp 1524952243
transform 1 0 1188 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1524952243
transform 1 0 1252 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1524952243
transform 1 0 1212 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1524952243
transform 1 0 1228 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1524952243
transform 1 0 1260 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2081
timestamp 1524952243
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1524952243
transform 1 0 1228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1524952243
transform 1 0 1236 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1524952243
transform 1 0 1188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1524952243
transform 1 0 1204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1524952243
transform 1 0 1220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1524952243
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1524952243
transform 1 0 1244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1524952243
transform 1 0 1260 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2438
timestamp 1524952243
transform 1 0 1188 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1524952243
transform 1 0 1220 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1524952243
transform 1 0 1260 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1524952243
transform 1 0 1276 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1524952243
transform 1 0 1268 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_2084
timestamp 1524952243
transform 1 0 1284 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2399
timestamp 1524952243
transform 1 0 1340 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2168
timestamp 1524952243
transform 1 0 1340 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2364
timestamp 1524952243
transform 1 0 1380 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1524952243
transform 1 0 1372 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2085
timestamp 1524952243
transform 1 0 1380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1524952243
transform 1 0 1364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1524952243
transform 1 0 1372 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2460
timestamp 1524952243
transform 1 0 1364 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1524952243
transform 1 0 1404 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1524952243
transform 1 0 1404 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2050
timestamp 1524952243
transform 1 0 1412 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1524952243
transform 1 0 1396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1524952243
transform 1 0 1396 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_2461
timestamp 1524952243
transform 1 0 1396 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1524952243
transform 1 0 1412 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1524952243
transform 1 0 1436 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1524952243
transform 1 0 1500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1524952243
transform 1 0 1444 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1524952243
transform 1 0 1468 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1524952243
transform 1 0 1508 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1524952243
transform 1 0 1444 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2087
timestamp 1524952243
transform 1 0 1436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1524952243
transform 1 0 1444 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2402
timestamp 1524952243
transform 1 0 1452 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2089
timestamp 1524952243
transform 1 0 1460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1524952243
transform 1 0 1468 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2403
timestamp 1524952243
transform 1 0 1476 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2091
timestamp 1524952243
transform 1 0 1524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1524952243
transform 1 0 1532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1524952243
transform 1 0 1428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1524952243
transform 1 0 1436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1524952243
transform 1 0 1452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1524952243
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1524952243
transform 1 0 1500 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2462
timestamp 1524952243
transform 1 0 1420 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_2093
timestamp 1524952243
transform 1 0 1580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1524952243
transform 1 0 1588 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2422
timestamp 1524952243
transform 1 0 1556 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2151
timestamp 1524952243
transform 1 0 1564 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2439
timestamp 1524952243
transform 1 0 1476 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1524952243
transform 1 0 1500 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1524952243
transform 1 0 1532 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1524952243
transform 1 0 1460 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1524952243
transform 1 0 1644 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1524952243
transform 1 0 1668 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2051
timestamp 1524952243
transform 1 0 1644 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_2394
timestamp 1524952243
transform 1 0 1652 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2095
timestamp 1524952243
transform 1 0 1636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1524952243
transform 1 0 1644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1524952243
transform 1 0 1652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1524952243
transform 1 0 1612 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2404
timestamp 1524952243
transform 1 0 1660 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1524952243
transform 1 0 1700 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2052
timestamp 1524952243
transform 1 0 1692 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1524952243
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1524952243
transform 1 0 1668 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1524952243
transform 1 0 1692 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_2154
timestamp 1524952243
transform 1 0 1700 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2442
timestamp 1524952243
transform 1 0 1676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1524952243
transform 1 0 1724 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1524952243
transform 1 0 1748 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2099
timestamp 1524952243
transform 1 0 1724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1524952243
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1524952243
transform 1 0 1756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1524952243
transform 1 0 1716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1524952243
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2423
timestamp 1524952243
transform 1 0 1748 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1524952243
transform 1 0 1740 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1524952243
transform 1 0 1764 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1524952243
transform 1 0 1812 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1524952243
transform 1 0 1780 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2102
timestamp 1524952243
transform 1 0 1780 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2396
timestamp 1524952243
transform 1 0 1836 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_2103
timestamp 1524952243
transform 1 0 1828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1524952243
transform 1 0 1836 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_2424
timestamp 1524952243
transform 1 0 1812 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1524952243
transform 1 0 1948 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1524952243
transform 1 0 1908 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_2105
timestamp 1524952243
transform 1 0 1892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1524952243
transform 1 0 1940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1524952243
transform 1 0 1836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1524952243
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2444
timestamp 1524952243
transform 1 0 1836 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1524952243
transform 1 0 1892 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_2159
timestamp 1524952243
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_2463
timestamp 1524952243
transform 1 0 1860 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1524952243
transform 1 0 1884 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1524952243
transform 1 0 1844 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1524952243
transform 1 0 1940 0 1 285
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_32
timestamp 1524952243
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_29
timestamp 1524952243
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_30
timestamp 1524952243
transform 1 0 80 0 -1 370
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_88
timestamp 1524952243
transform -1 0 184 0 -1 370
box -8 -3 104 105
use FILL  FILL_31
timestamp 1524952243
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_32
timestamp 1524952243
transform 1 0 192 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_80
timestamp 1524952243
transform -1 0 232 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1524952243
transform -1 0 264 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1524952243
transform -1 0 296 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1524952243
transform -1 0 328 0 -1 370
box -8 -3 34 105
use M3_M2  M3_M2_2486
timestamp 1524952243
transform 1 0 356 0 1 275
box -3 -3 3 3
use NOR2X1  NOR2X1_46
timestamp 1524952243
transform 1 0 328 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_128
timestamp 1524952243
transform 1 0 352 0 -1 370
box -9 -3 26 105
use XNOR2X1  XNOR2X1_54
timestamp 1524952243
transform -1 0 424 0 -1 370
box -8 -3 64 105
use AND2X2  AND2X2_23
timestamp 1524952243
transform -1 0 456 0 -1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_84
timestamp 1524952243
transform -1 0 488 0 -1 370
box -8 -3 34 105
use NAND3X1  NAND3X1_26
timestamp 1524952243
transform 1 0 488 0 -1 370
box -8 -3 40 105
use FILL  FILL_33
timestamp 1524952243
transform 1 0 520 0 -1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_55
timestamp 1524952243
transform -1 0 584 0 -1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_55
timestamp 1524952243
transform 1 0 584 0 -1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_56
timestamp 1524952243
transform 1 0 640 0 -1 370
box -8 -3 64 105
use NOR2X1  NOR2X1_47
timestamp 1524952243
transform 1 0 696 0 -1 370
box -8 -3 32 105
use XOR2X1  XOR2X1_56
timestamp 1524952243
transform 1 0 720 0 -1 370
box -8 -3 64 105
use FILL  FILL_34
timestamp 1524952243
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_35
timestamp 1524952243
transform 1 0 784 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_75
timestamp 1524952243
transform 1 0 792 0 -1 370
box -8 -3 46 105
use AND2X2  AND2X2_24
timestamp 1524952243
transform 1 0 832 0 -1 370
box -8 -3 40 105
use FILL  FILL_36
timestamp 1524952243
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_37
timestamp 1524952243
transform 1 0 872 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_2487
timestamp 1524952243
transform 1 0 892 0 1 275
box -3 -3 3 3
use FILL  FILL_38
timestamp 1524952243
transform 1 0 880 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_2488
timestamp 1524952243
transform 1 0 908 0 1 275
box -3 -3 3 3
use FILL  FILL_39
timestamp 1524952243
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_40
timestamp 1524952243
transform 1 0 896 0 -1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_57
timestamp 1524952243
transform 1 0 904 0 -1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_57
timestamp 1524952243
transform -1 0 1016 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_58
timestamp 1524952243
transform 1 0 1016 0 -1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_58
timestamp 1524952243
transform 1 0 1072 0 -1 370
box -8 -3 64 105
use FILL  FILL_41
timestamp 1524952243
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_42
timestamp 1524952243
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_43
timestamp 1524952243
transform 1 0 1144 0 -1 370
box -8 -3 32 105
use FILL  FILL_43
timestamp 1524952243
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_2489
timestamp 1524952243
transform 1 0 1188 0 1 275
box -3 -3 3 3
use FILL  FILL_44
timestamp 1524952243
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_76
timestamp 1524952243
transform -1 0 1224 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_2490
timestamp 1524952243
transform 1 0 1236 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_77
timestamp 1524952243
transform 1 0 1224 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_2491
timestamp 1524952243
transform 1 0 1284 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1524952243
transform 1 0 1300 0 1 275
box -3 -3 3 3
use FILL  FILL_45
timestamp 1524952243
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_46
timestamp 1524952243
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_59
timestamp 1524952243
transform -1 0 1336 0 -1 370
box -8 -3 64 105
use FILL  FILL_47
timestamp 1524952243
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_85
timestamp 1524952243
transform -1 0 1376 0 -1 370
box -8 -3 34 105
use NAND2X1  NAND2X1_44
timestamp 1524952243
transform 1 0 1376 0 -1 370
box -8 -3 32 105
use FILL  FILL_48
timestamp 1524952243
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_48
timestamp 1524952243
transform 1 0 1408 0 -1 370
box -8 -3 32 105
use AOI22X1  AOI22X1_78
timestamp 1524952243
transform -1 0 1472 0 -1 370
box -8 -3 46 105
use XOR2X1  XOR2X1_59
timestamp 1524952243
transform 1 0 1472 0 -1 370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_60
timestamp 1524952243
transform 1 0 1528 0 -1 370
box -8 -3 64 105
use M3_M2  M3_M2_2493
timestamp 1524952243
transform 1 0 1620 0 1 275
box -3 -3 3 3
use XOR2X1  XOR2X1_60
timestamp 1524952243
transform 1 0 1584 0 -1 370
box -8 -3 64 105
use NOR2X1  NOR2X1_49
timestamp 1524952243
transform 1 0 1640 0 -1 370
box -8 -3 32 105
use AOI21X1  AOI21X1_10
timestamp 1524952243
transform 1 0 1664 0 -1 370
box -7 -3 39 105
use INVX2  INVX2_129
timestamp 1524952243
transform 1 0 1696 0 -1 370
box -9 -3 26 105
use FILL  FILL_49
timestamp 1524952243
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_79
timestamp 1524952243
transform -1 0 1760 0 -1 370
box -8 -3 46 105
use FILL  FILL_50
timestamp 1524952243
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_51
timestamp 1524952243
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_61
timestamp 1524952243
transform 1 0 1776 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_61
timestamp 1524952243
transform 1 0 1832 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_62
timestamp 1524952243
transform -1 0 1944 0 -1 370
box -8 -3 64 105
use top_module_VIA0  top_module_VIA0_33
timestamp 1524952243
transform 1 0 1994 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_2520
timestamp 1524952243
transform 1 0 76 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2206
timestamp 1524952243
transform 1 0 76 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1524952243
transform 1 0 196 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1524952243
transform 1 0 156 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1524952243
transform 1 0 196 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1524952243
transform 1 0 228 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2182
timestamp 1524952243
transform 1 0 228 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1524952243
transform 1 0 220 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2566
timestamp 1524952243
transform 1 0 228 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2280
timestamp 1524952243
transform 1 0 180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1524952243
transform 1 0 196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1524952243
transform 1 0 220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1524952243
transform 1 0 228 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2606
timestamp 1524952243
transform 1 0 156 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1524952243
transform 1 0 196 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1524952243
transform 1 0 228 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1524952243
transform 1 0 220 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_2209
timestamp 1524952243
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1524952243
transform 1 0 260 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_2516
timestamp 1524952243
transform 1 0 316 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1524952243
transform 1 0 292 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1524952243
transform 1 0 276 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2284
timestamp 1524952243
transform 1 0 284 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2625
timestamp 1524952243
transform 1 0 284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1524952243
transform 1 0 340 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2210
timestamp 1524952243
transform 1 0 292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1524952243
transform 1 0 300 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2568
timestamp 1524952243
transform 1 0 308 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1524952243
transform 1 0 396 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1524952243
transform 1 0 380 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2212
timestamp 1524952243
transform 1 0 316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1524952243
transform 1 0 332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1524952243
transform 1 0 340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1524952243
transform 1 0 356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1524952243
transform 1 0 300 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2592
timestamp 1524952243
transform 1 0 316 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1524952243
transform 1 0 364 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1524952243
transform 1 0 460 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1524952243
transform 1 0 436 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1524952243
transform 1 0 476 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1524952243
transform 1 0 476 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1524952243
transform 1 0 444 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2216
timestamp 1524952243
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1524952243
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1524952243
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1524952243
transform 1 0 444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1524952243
transform 1 0 452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1524952243
transform 1 0 324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1524952243
transform 1 0 332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1524952243
transform 1 0 364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1524952243
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1524952243
transform 1 0 388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1524952243
transform 1 0 404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1524952243
transform 1 0 412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2626
timestamp 1524952243
transform 1 0 324 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1524952243
transform 1 0 372 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_2221
timestamp 1524952243
transform 1 0 484 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2570
timestamp 1524952243
transform 1 0 492 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2293
timestamp 1524952243
transform 1 0 476 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2628
timestamp 1524952243
transform 1 0 412 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1524952243
transform 1 0 460 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1524952243
transform 1 0 580 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1524952243
transform 1 0 604 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1524952243
transform 1 0 620 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1524952243
transform 1 0 636 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_2171
timestamp 1524952243
transform 1 0 540 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1524952243
transform 1 0 556 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1524952243
transform 1 0 508 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1524952243
transform 1 0 524 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1524952243
transform 1 0 500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2609
timestamp 1524952243
transform 1 0 500 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1524952243
transform 1 0 540 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2185
timestamp 1524952243
transform 1 0 556 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2537
timestamp 1524952243
transform 1 0 564 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1524952243
transform 1 0 612 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2222
timestamp 1524952243
transform 1 0 524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1524952243
transform 1 0 548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1524952243
transform 1 0 524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2593
timestamp 1524952243
transform 1 0 532 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1524952243
transform 1 0 484 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1524952243
transform 1 0 508 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1524952243
transform 1 0 556 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2224
timestamp 1524952243
transform 1 0 564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1524952243
transform 1 0 580 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2572
timestamp 1524952243
transform 1 0 588 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1524952243
transform 1 0 668 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1524952243
transform 1 0 652 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2226
timestamp 1524952243
transform 1 0 612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1524952243
transform 1 0 636 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2573
timestamp 1524952243
transform 1 0 644 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1524952243
transform 1 0 668 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2186
timestamp 1524952243
transform 1 0 676 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1524952243
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1524952243
transform 1 0 668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1524952243
transform 1 0 628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2594
timestamp 1524952243
transform 1 0 636 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2297
timestamp 1524952243
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1524952243
transform 1 0 660 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2632
timestamp 1524952243
transform 1 0 588 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1524952243
transform 1 0 620 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1524952243
transform 1 0 676 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2173
timestamp 1524952243
transform 1 0 724 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_2540
timestamp 1524952243
transform 1 0 732 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1524952243
transform 1 0 780 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_2187
timestamp 1524952243
transform 1 0 740 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2541
timestamp 1524952243
transform 1 0 764 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1524952243
transform 1 0 788 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_2188
timestamp 1524952243
transform 1 0 772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1524952243
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1524952243
transform 1 0 732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1524952243
transform 1 0 676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2595
timestamp 1524952243
transform 1 0 692 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1524952243
transform 1 0 676 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1524952243
transform 1 0 676 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1524952243
transform 1 0 740 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2232
timestamp 1524952243
transform 1 0 748 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2596
timestamp 1524952243
transform 1 0 732 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2300
timestamp 1524952243
transform 1 0 748 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2611
timestamp 1524952243
transform 1 0 748 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1524952243
transform 1 0 724 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1524952243
transform 1 0 748 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1524952243
transform 1 0 780 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1524952243
transform 1 0 844 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1524952243
transform 1 0 828 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1524952243
transform 1 0 820 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1524952243
transform 1 0 852 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1524952243
transform 1 0 868 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1524952243
transform 1 0 900 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1524952243
transform 1 0 908 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1524952243
transform 1 0 892 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2545
timestamp 1524952243
transform 1 0 900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1524952243
transform 1 0 972 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1524952243
transform 1 0 948 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2190
timestamp 1524952243
transform 1 0 916 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1524952243
transform 1 0 788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1524952243
transform 1 0 804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1524952243
transform 1 0 828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1524952243
transform 1 0 844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1524952243
transform 1 0 852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1524952243
transform 1 0 868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1524952243
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1524952243
transform 1 0 772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1524952243
transform 1 0 780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2597
timestamp 1524952243
transform 1 0 788 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2303
timestamp 1524952243
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1524952243
transform 1 0 820 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2612
timestamp 1524952243
transform 1 0 796 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1524952243
transform 1 0 828 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1524952243
transform 1 0 892 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1524952243
transform 1 0 932 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1524952243
transform 1 0 956 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2240
timestamp 1524952243
transform 1 0 900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1524952243
transform 1 0 852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1524952243
transform 1 0 860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1524952243
transform 1 0 876 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1524952243
transform 1 0 884 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1524952243
transform 1 0 852 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1524952243
transform 1 0 836 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1524952243
transform 1 0 876 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1524952243
transform 1 0 892 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1524952243
transform 1 0 924 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2241
timestamp 1524952243
transform 1 0 932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1524952243
transform 1 0 924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1524952243
transform 1 0 1012 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1524952243
transform 1 0 1028 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_2548
timestamp 1524952243
transform 1 0 1004 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2191
timestamp 1524952243
transform 1 0 1012 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2549
timestamp 1524952243
transform 1 0 1020 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2242
timestamp 1524952243
transform 1 0 972 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1524952243
transform 1 0 1012 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1524952243
transform 1 0 1060 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2192
timestamp 1524952243
transform 1 0 1076 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1524952243
transform 1 0 1020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1524952243
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1524952243
transform 1 0 1004 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1524952243
transform 1 0 1004 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1524952243
transform 1 0 972 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1524952243
transform 1 0 988 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1524952243
transform 1 0 1052 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1524952243
transform 1 0 1100 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2193
timestamp 1524952243
transform 1 0 1108 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1524952243
transform 1 0 1076 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1524952243
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1524952243
transform 1 0 1100 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2600
timestamp 1524952243
transform 1 0 1060 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2310
timestamp 1524952243
transform 1 0 1068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1524952243
transform 1 0 1076 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2601
timestamp 1524952243
transform 1 0 1092 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2312
timestamp 1524952243
transform 1 0 1100 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2615
timestamp 1524952243
transform 1 0 1076 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1524952243
transform 1 0 1140 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1524952243
transform 1 0 1124 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2177
timestamp 1524952243
transform 1 0 1140 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1524952243
transform 1 0 1124 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1524952243
transform 1 0 1156 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2552
timestamp 1524952243
transform 1 0 1164 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2248
timestamp 1524952243
transform 1 0 1148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1524952243
transform 1 0 1124 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2616
timestamp 1524952243
transform 1 0 1124 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1524952243
transform 1 0 1156 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2249
timestamp 1524952243
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1524952243
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1524952243
transform 1 0 1172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2602
timestamp 1524952243
transform 1 0 1180 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1524952243
transform 1 0 1164 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1524952243
transform 1 0 1204 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1524952243
transform 1 0 1196 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_2178
timestamp 1524952243
transform 1 0 1244 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1524952243
transform 1 0 1228 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1524952243
transform 1 0 1188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1524952243
transform 1 0 1212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1524952243
transform 1 0 1188 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2553
timestamp 1524952243
transform 1 0 1236 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1524952243
transform 1 0 1276 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_2197
timestamp 1524952243
transform 1 0 1252 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2554
timestamp 1524952243
transform 1 0 1276 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1524952243
transform 1 0 1348 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1524952243
transform 1 0 1332 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1524952243
transform 1 0 1340 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1524952243
transform 1 0 1364 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2253
timestamp 1524952243
transform 1 0 1236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1524952243
transform 1 0 1260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1524952243
transform 1 0 1276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1524952243
transform 1 0 1292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1524952243
transform 1 0 1300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1524952243
transform 1 0 1220 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1524952243
transform 1 0 1204 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1524952243
transform 1 0 1260 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1524952243
transform 1 0 1308 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2258
timestamp 1524952243
transform 1 0 1316 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2583
timestamp 1524952243
transform 1 0 1332 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1524952243
transform 1 0 1460 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1524952243
transform 1 0 1452 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1524952243
transform 1 0 1420 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1524952243
transform 1 0 1444 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2198
timestamp 1524952243
transform 1 0 1452 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1524952243
transform 1 0 1340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1524952243
transform 1 0 1364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1524952243
transform 1 0 1388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1524952243
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1524952243
transform 1 0 1268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1524952243
transform 1 0 1300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1524952243
transform 1 0 1308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2604
timestamp 1524952243
transform 1 0 1316 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2320
timestamp 1524952243
transform 1 0 1324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1524952243
transform 1 0 1340 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1524952243
transform 1 0 1428 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2263
timestamp 1524952243
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1524952243
transform 1 0 1396 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2617
timestamp 1524952243
transform 1 0 1292 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1524952243
transform 1 0 1324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1524952243
transform 1 0 1340 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1524952243
transform 1 0 1284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1524952243
transform 1 0 1484 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2264
timestamp 1524952243
transform 1 0 1468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1524952243
transform 1 0 1452 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2620
timestamp 1524952243
transform 1 0 1452 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_2324
timestamp 1524952243
transform 1 0 1476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1524952243
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2559
timestamp 1524952243
transform 1 0 1556 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2265
timestamp 1524952243
transform 1 0 1532 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2585
timestamp 1524952243
transform 1 0 1540 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1524952243
transform 1 0 1612 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2199
timestamp 1524952243
transform 1 0 1652 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1524952243
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1524952243
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1524952243
transform 1 0 1620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1524952243
transform 1 0 1644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1524952243
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1524952243
transform 1 0 1596 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2621
timestamp 1524952243
transform 1 0 1596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1524952243
transform 1 0 1676 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1524952243
transform 1 0 1660 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2270
timestamp 1524952243
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1524952243
transform 1 0 1676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1524952243
transform 1 0 1652 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1524952243
transform 1 0 1676 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_2329
timestamp 1524952243
transform 1 0 1684 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2645
timestamp 1524952243
transform 1 0 1668 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1524952243
transform 1 0 1708 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1524952243
transform 1 0 1748 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1524952243
transform 1 0 1740 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_2200
timestamp 1524952243
transform 1 0 1700 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2561
timestamp 1524952243
transform 1 0 1724 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2201
timestamp 1524952243
transform 1 0 1732 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2587
timestamp 1524952243
transform 1 0 1700 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2330
timestamp 1524952243
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2514
timestamp 1524952243
transform 1 0 1820 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1524952243
transform 1 0 1796 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2272
timestamp 1524952243
transform 1 0 1740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1524952243
transform 1 0 1756 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_2588
timestamp 1524952243
transform 1 0 1764 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1524952243
transform 1 0 1788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1524952243
transform 1 0 1796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1524952243
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1524952243
transform 1 0 1732 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2622
timestamp 1524952243
transform 1 0 1732 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_2332
timestamp 1524952243
transform 1 0 1788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1524952243
transform 1 0 1796 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2646
timestamp 1524952243
transform 1 0 1748 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1524952243
transform 1 0 1860 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_2202
timestamp 1524952243
transform 1 0 1868 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2563
timestamp 1524952243
transform 1 0 1876 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1524952243
transform 1 0 1860 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1524952243
transform 1 0 1916 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_2179
timestamp 1524952243
transform 1 0 1916 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1524952243
transform 1 0 1924 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1524952243
transform 1 0 1900 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1524952243
transform 1 0 1908 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1524952243
transform 1 0 1916 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_2205
timestamp 1524952243
transform 1 0 1932 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1524952243
transform 1 0 1876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1524952243
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1524952243
transform 1 0 1844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1524952243
transform 1 0 1852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1524952243
transform 1 0 1868 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1524952243
transform 1 0 1860 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1524952243
transform 1 0 1812 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1524952243
transform 1 0 1844 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1524952243
transform 1 0 1900 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_2279
timestamp 1524952243
transform 1 0 1916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1524952243
transform 1 0 1900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_2591
timestamp 1524952243
transform 1 0 1932 0 1 215
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_34
timestamp 1524952243
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_52
timestamp 1524952243
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_54
timestamp 1524952243
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_56
timestamp 1524952243
transform 1 0 88 0 1 170
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_89
timestamp 1524952243
transform -1 0 192 0 1 170
box -8 -3 104 105
use OAI21X1  OAI21X1_86
timestamp 1524952243
transform -1 0 224 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1524952243
transform -1 0 256 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_50
timestamp 1524952243
transform 1 0 256 0 1 170
box -8 -3 32 105
use INVX2  INVX2_130
timestamp 1524952243
transform 1 0 280 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_80
timestamp 1524952243
transform -1 0 336 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1524952243
transform 1 0 336 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1524952243
transform -1 0 416 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_2649
timestamp 1524952243
transform 1 0 468 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_63
timestamp 1524952243
transform 1 0 416 0 1 170
box -8 -3 64 105
use OAI21X1  OAI21X1_88
timestamp 1524952243
transform 1 0 472 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_45
timestamp 1524952243
transform -1 0 528 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_27
timestamp 1524952243
transform -1 0 560 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_2650
timestamp 1524952243
transform 1 0 580 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_64
timestamp 1524952243
transform -1 0 616 0 1 170
box -8 -3 64 105
use AOI22X1  AOI22X1_83
timestamp 1524952243
transform -1 0 656 0 1 170
box -8 -3 46 105
use NAND2X1  NAND2X1_46
timestamp 1524952243
transform 1 0 656 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_89
timestamp 1524952243
transform 1 0 680 0 1 170
box -8 -3 34 105
use NAND3X1  NAND3X1_28
timestamp 1524952243
transform -1 0 744 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_2651
timestamp 1524952243
transform 1 0 756 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_90
timestamp 1524952243
transform 1 0 744 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_2652
timestamp 1524952243
transform 1 0 804 0 1 175
box -3 -3 3 3
use AND2X2  AND2X2_25
timestamp 1524952243
transform 1 0 776 0 1 170
box -8 -3 40 105
use AOI22X1  AOI22X1_84
timestamp 1524952243
transform 1 0 808 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1524952243
transform -1 0 888 0 1 170
box -8 -3 46 105
use NAND3X1  NAND3X1_29
timestamp 1524952243
transform 1 0 888 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1524952243
transform 1 0 920 0 1 170
box -8 -3 40 105
use XNOR2X1  XNOR2X1_62
timestamp 1524952243
transform -1 0 1008 0 1 170
box -8 -3 64 105
use NAND3X1  NAND3X1_30
timestamp 1524952243
transform 1 0 1008 0 1 170
box -8 -3 40 105
use OAI21X1  OAI21X1_91
timestamp 1524952243
transform -1 0 1072 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1524952243
transform -1 0 1104 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_47
timestamp 1524952243
transform -1 0 1128 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_31
timestamp 1524952243
transform -1 0 1160 0 1 170
box -8 -3 40 105
use INVX2  INVX2_131
timestamp 1524952243
transform -1 0 1176 0 1 170
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1524952243
transform -1 0 1192 0 1 170
box -9 -3 26 105
use AND2X2  AND2X2_27
timestamp 1524952243
transform -1 0 1224 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_2653
timestamp 1524952243
transform 1 0 1244 0 1 175
box -3 -3 3 3
use NAND3X1  NAND3X1_32
timestamp 1524952243
transform 1 0 1224 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_2654
timestamp 1524952243
transform 1 0 1268 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1524952243
transform 1 0 1316 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_86
timestamp 1524952243
transform 1 0 1256 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_2656
timestamp 1524952243
transform 1 0 1332 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_87
timestamp 1524952243
transform 1 0 1296 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_2657
timestamp 1524952243
transform 1 0 1380 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_65
timestamp 1524952243
transform 1 0 1336 0 1 170
box -8 -3 64 105
use M3_M2  M3_M2_2658
timestamp 1524952243
transform 1 0 1436 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_66
timestamp 1524952243
transform 1 0 1392 0 1 170
box -8 -3 64 105
use M3_M2  M3_M2_2659
timestamp 1524952243
transform 1 0 1460 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1524952243
transform 1 0 1476 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_93
timestamp 1524952243
transform -1 0 1480 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_2661
timestamp 1524952243
transform 1 0 1524 0 1 175
box -3 -3 3 3
use XNOR2X1  XNOR2X1_63
timestamp 1524952243
transform -1 0 1536 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_64
timestamp 1524952243
transform -1 0 1592 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_67
timestamp 1524952243
transform 1 0 1592 0 1 170
box -8 -3 64 105
use OAI21X1  OAI21X1_94
timestamp 1524952243
transform -1 0 1680 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_2662
timestamp 1524952243
transform 1 0 1708 0 1 175
box -3 -3 3 3
use NAND2X1  NAND2X1_48
timestamp 1524952243
transform 1 0 1680 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_2663
timestamp 1524952243
transform 1 0 1732 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_95
timestamp 1524952243
transform 1 0 1704 0 1 170
box -8 -3 34 105
use XNOR2X1  XNOR2X1_65
timestamp 1524952243
transform -1 0 1792 0 1 170
box -8 -3 64 105
use M3_M2  M3_M2_2664
timestamp 1524952243
transform 1 0 1820 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1524952243
transform 1 0 1852 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_68
timestamp 1524952243
transform -1 0 1848 0 1 170
box -8 -3 64 105
use NAND2X1  NAND2X1_49
timestamp 1524952243
transform 1 0 1848 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_96
timestamp 1524952243
transform 1 0 1872 0 1 170
box -8 -3 34 105
use NAND3X1  NAND3X1_33
timestamp 1524952243
transform 1 0 1904 0 1 170
box -8 -3 40 105
use FILL  FILL_57
timestamp 1524952243
transform 1 0 1936 0 1 170
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_35
timestamp 1524952243
transform 1 0 1970 0 1 170
box -10 -3 10 3
use top_module_VIA0  top_module_VIA0_36
timestamp 1524952243
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_53
timestamp 1524952243
transform 1 0 72 0 -1 170
box -8 -3 16 105
use FILL  FILL_55
timestamp 1524952243
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_58
timestamp 1524952243
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_59
timestamp 1524952243
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_60
timestamp 1524952243
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_61
timestamp 1524952243
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_62
timestamp 1524952243
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_63
timestamp 1524952243
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_64
timestamp 1524952243
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_65
timestamp 1524952243
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_66
timestamp 1524952243
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_67
timestamp 1524952243
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_68
timestamp 1524952243
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_69
timestamp 1524952243
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_70
timestamp 1524952243
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_71
timestamp 1524952243
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_72
timestamp 1524952243
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_73
timestamp 1524952243
transform 1 0 208 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_2341
timestamp 1524952243
transform 1 0 228 0 1 135
box -2 -2 2 2
use FILL  FILL_74
timestamp 1524952243
transform 1 0 216 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_2384
timestamp 1524952243
transform 1 0 260 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2688
timestamp 1524952243
transform 1 0 292 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1524952243
transform 1 0 332 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1524952243
transform 1 0 348 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2342
timestamp 1524952243
transform 1 0 308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1524952243
transform 1 0 316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1524952243
transform 1 0 300 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2737
timestamp 1524952243
transform 1 0 260 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1524952243
transform 1 0 276 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1524952243
transform 1 0 292 0 1 115
box -3 -3 3 3
use XNOR2X1  XNOR2X1_66
timestamp 1524952243
transform 1 0 224 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2666
timestamp 1524952243
transform 1 0 388 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1524952243
transform 1 0 372 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1524952243
transform 1 0 436 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1524952243
transform 1 0 452 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1524952243
transform 1 0 428 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2344
timestamp 1524952243
transform 1 0 372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1524952243
transform 1 0 420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1524952243
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1524952243
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1524952243
transform 1 0 364 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2740
timestamp 1524952243
transform 1 0 340 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1524952243
transform 1 0 308 0 1 105
box -3 -3 3 3
use AND2X2  AND2X2_28
timestamp 1524952243
transform -1 0 312 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_2722
timestamp 1524952243
transform 1 0 420 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2388
timestamp 1524952243
transform 1 0 428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1524952243
transform 1 0 428 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_2761
timestamp 1524952243
transform 1 0 364 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1524952243
transform 1 0 412 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1524952243
transform 1 0 428 0 1 105
box -3 -3 3 3
use XOR2X1  XOR2X1_69
timestamp 1524952243
transform 1 0 312 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2778
timestamp 1524952243
transform 1 0 428 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_70
timestamp 1524952243
transform 1 0 368 0 -1 170
box -8 -3 64 105
use M2_M1  M2_M1_2347
timestamp 1524952243
transform 1 0 452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1524952243
transform 1 0 460 0 1 125
box -2 -2 2 2
use OAI21X1  OAI21X1_97
timestamp 1524952243
transform -1 0 456 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_2669
timestamp 1524952243
transform 1 0 476 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_2339
timestamp 1524952243
transform 1 0 476 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_2723
timestamp 1524952243
transform 1 0 476 0 1 125
box -3 -3 3 3
use INVX2  INVX2_133
timestamp 1524952243
transform -1 0 472 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_2700
timestamp 1524952243
transform 1 0 500 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1524952243
transform 1 0 508 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1524952243
transform 1 0 500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1524952243
transform 1 0 508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1524952243
transform 1 0 500 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2724
timestamp 1524952243
transform 1 0 508 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1524952243
transform 1 0 492 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1524952243
transform 1 0 524 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1524952243
transform 1 0 524 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1524952243
transform 1 0 612 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1524952243
transform 1 0 684 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2350
timestamp 1524952243
transform 1 0 580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1524952243
transform 1 0 596 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2713
timestamp 1524952243
transform 1 0 604 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2352
timestamp 1524952243
transform 1 0 612 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2714
timestamp 1524952243
transform 1 0 628 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2353
timestamp 1524952243
transform 1 0 676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1524952243
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1524952243
transform 1 0 524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1524952243
transform 1 0 532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1524952243
transform 1 0 548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1524952243
transform 1 0 580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1524952243
transform 1 0 604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1524952243
transform 1 0 620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1524952243
transform 1 0 628 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2741
timestamp 1524952243
transform 1 0 532 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1524952243
transform 1 0 516 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1524952243
transform 1 0 500 0 1 85
box -3 -3 3 3
use AOI21X1  AOI21X1_11
timestamp 1524952243
transform -1 0 504 0 -1 170
box -7 -3 39 105
use NOR2X1  NOR2X1_51
timestamp 1524952243
transform 1 0 504 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_2742
timestamp 1524952243
transform 1 0 580 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1524952243
transform 1 0 548 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1524952243
transform 1 0 588 0 1 85
box -3 -3 3 3
use XOR2X1  XOR2X1_71
timestamp 1524952243
transform -1 0 584 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2743
timestamp 1524952243
transform 1 0 628 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1524952243
transform 1 0 620 0 1 105
box -3 -3 3 3
use AOI22X1  AOI22X1_88
timestamp 1524952243
transform 1 0 584 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_2793
timestamp 1524952243
transform 1 0 684 0 1 75
box -3 -3 3 3
use XNOR2X1  XNOR2X1_67
timestamp 1524952243
transform -1 0 680 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2671
timestamp 1524952243
transform 1 0 740 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_2355
timestamp 1524952243
transform 1 0 732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1524952243
transform 1 0 740 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2715
timestamp 1524952243
transform 1 0 764 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2357
timestamp 1524952243
transform 1 0 772 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2672
timestamp 1524952243
transform 1 0 828 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1524952243
transform 1 0 860 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1524952243
transform 1 0 884 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1524952243
transform 1 0 820 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2358
timestamp 1524952243
transform 1 0 828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1524952243
transform 1 0 732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1524952243
transform 1 0 748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1524952243
transform 1 0 772 0 1 125
box -2 -2 2 2
use XOR2X1  XOR2X1_72
timestamp 1524952243
transform 1 0 680 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2725
timestamp 1524952243
transform 1 0 796 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1524952243
transform 1 0 884 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2359
timestamp 1524952243
transform 1 0 876 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2705
timestamp 1524952243
transform 1 0 948 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1524952243
transform 1 0 980 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2360
timestamp 1524952243
transform 1 0 940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1524952243
transform 1 0 948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1524952243
transform 1 0 804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1524952243
transform 1 0 820 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1524952243
transform 1 0 852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1524952243
transform 1 0 884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1524952243
transform 1 0 908 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2744
timestamp 1524952243
transform 1 0 772 0 1 115
box -3 -3 3 3
use AND2X2  AND2X2_29
timestamp 1524952243
transform 1 0 736 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_2745
timestamp 1524952243
transform 1 0 820 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1524952243
transform 1 0 852 0 1 115
box -3 -3 3 3
use XNOR2X1  XNOR2X1_68
timestamp 1524952243
transform 1 0 768 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2766
timestamp 1524952243
transform 1 0 908 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1524952243
transform 1 0 884 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_73
timestamp 1524952243
transform 1 0 824 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_74
timestamp 1524952243
transform 1 0 880 0 -1 170
box -8 -3 64 105
use M2_M1  M2_M1_2406
timestamp 1524952243
transform 1 0 956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1524952243
transform 1 0 972 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1524952243
transform 1 0 980 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2747
timestamp 1524952243
transform 1 0 980 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1524952243
transform 1 0 956 0 1 85
box -3 -3 3 3
use AOI22X1  AOI22X1_89
timestamp 1524952243
transform -1 0 976 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_2707
timestamp 1524952243
transform 1 0 1036 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1524952243
transform 1 0 1076 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1524952243
transform 1 0 1068 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2362
timestamp 1524952243
transform 1 0 1036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1524952243
transform 1 0 1044 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1524952243
transform 1 0 1060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1524952243
transform 1 0 1076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1524952243
transform 1 0 1028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1524952243
transform 1 0 1036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1524952243
transform 1 0 1052 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1524952243
transform 1 0 1068 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2748
timestamp 1524952243
transform 1 0 1060 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1524952243
transform 1 0 1036 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_75
timestamp 1524952243
transform 1 0 976 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2794
timestamp 1524952243
transform 1 0 1044 0 1 75
box -3 -3 3 3
use AOI22X1  AOI22X1_90
timestamp 1524952243
transform 1 0 1032 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_2676
timestamp 1524952243
transform 1 0 1172 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1524952243
transform 1 0 1124 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1524952243
transform 1 0 1212 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1524952243
transform 1 0 1204 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2366
timestamp 1524952243
transform 1 0 1180 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1524952243
transform 1 0 1188 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1524952243
transform 1 0 1244 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_2367
timestamp 1524952243
transform 1 0 1196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1524952243
transform 1 0 1212 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1524952243
transform 1 0 1124 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1524952243
transform 1 0 1132 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2726
timestamp 1524952243
transform 1 0 1148 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1524952243
transform 1 0 1220 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2415
timestamp 1524952243
transform 1 0 1180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1524952243
transform 1 0 1188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1524952243
transform 1 0 1204 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1524952243
transform 1 0 1132 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1524952243
transform 1 0 1100 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1524952243
transform 1 0 1124 0 1 75
box -3 -3 3 3
use XNOR2X1  XNOR2X1_69
timestamp 1524952243
transform -1 0 1128 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2727
timestamp 1524952243
transform 1 0 1212 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1524952243
transform 1 0 1300 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1524952243
transform 1 0 1292 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2369
timestamp 1524952243
transform 1 0 1276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1524952243
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2720
timestamp 1524952243
transform 1 0 1300 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2371
timestamp 1524952243
transform 1 0 1308 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2721
timestamp 1524952243
transform 1 0 1316 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_2372
timestamp 1524952243
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1524952243
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1524952243
transform 1 0 1252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1524952243
transform 1 0 1284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1524952243
transform 1 0 1300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1524952243
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1524952243
transform 1 0 1324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1524952243
transform 1 0 1348 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2749
timestamp 1524952243
transform 1 0 1180 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1524952243
transform 1 0 1188 0 1 105
box -3 -3 3 3
use XNOR2X1  XNOR2X1_70
timestamp 1524952243
transform 1 0 1128 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2750
timestamp 1524952243
transform 1 0 1220 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1524952243
transform 1 0 1196 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1524952243
transform 1 0 1212 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1524952243
transform 1 0 1204 0 1 85
box -3 -3 3 3
use AOI22X1  AOI22X1_91
timestamp 1524952243
transform 1 0 1184 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_2751
timestamp 1524952243
transform 1 0 1284 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1524952243
transform 1 0 1252 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1524952243
transform 1 0 1268 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1524952243
transform 1 0 1268 0 1 75
box -3 -3 3 3
use XOR2X1  XOR2X1_76
timestamp 1524952243
transform -1 0 1280 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2728
timestamp 1524952243
transform 1 0 1380 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1524952243
transform 1 0 1428 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1524952243
transform 1 0 1468 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2373
timestamp 1524952243
transform 1 0 1444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1524952243
transform 1 0 1388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1524952243
transform 1 0 1404 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2752
timestamp 1524952243
transform 1 0 1348 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1524952243
transform 1 0 1324 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1524952243
transform 1 0 1316 0 1 95
box -3 -3 3 3
use AOI22X1  AOI22X1_92
timestamp 1524952243
transform 1 0 1280 0 -1 170
box -8 -3 46 105
use XOR2X1  XOR2X1_77
timestamp 1524952243
transform 1 0 1320 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2729
timestamp 1524952243
transform 1 0 1412 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2427
timestamp 1524952243
transform 1 0 1420 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2730
timestamp 1524952243
transform 1 0 1428 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1524952243
transform 1 0 1404 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_2449
timestamp 1524952243
transform 1 0 1412 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1524952243
transform 1 0 1460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1524952243
transform 1 0 1436 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_2754
timestamp 1524952243
transform 1 0 1444 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1524952243
transform 1 0 1460 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1524952243
transform 1 0 1516 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2374
timestamp 1524952243
transform 1 0 1532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1524952243
transform 1 0 1516 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1524952243
transform 1 0 1524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1524952243
transform 1 0 1532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1524952243
transform 1 0 1500 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_2771
timestamp 1524952243
transform 1 0 1388 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1524952243
transform 1 0 1404 0 1 105
box -3 -3 3 3
use M2_M1  M2_M1_2456
timestamp 1524952243
transform 1 0 1412 0 1 105
box -2 -2 2 2
use M3_M2  M3_M2_2773
timestamp 1524952243
transform 1 0 1420 0 1 105
box -3 -3 3 3
use AND2X2  AND2X2_30
timestamp 1524952243
transform 1 0 1376 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1524952243
transform 1 0 1408 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_2774
timestamp 1524952243
transform 1 0 1500 0 1 105
box -3 -3 3 3
use XNOR2X1  XNOR2X1_71
timestamp 1524952243
transform -1 0 1496 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2775
timestamp 1524952243
transform 1 0 1532 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1524952243
transform 1 0 1524 0 1 85
box -3 -3 3 3
use OAI21X1  OAI21X1_98
timestamp 1524952243
transform -1 0 1528 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_2694
timestamp 1524952243
transform 1 0 1548 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1524952243
transform 1 0 1604 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1524952243
transform 1 0 1652 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_2375
timestamp 1524952243
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1524952243
transform 1 0 1556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1524952243
transform 1 0 1572 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2731
timestamp 1524952243
transform 1 0 1580 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2376
timestamp 1524952243
transform 1 0 1660 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1524952243
transform 1 0 1612 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1524952243
transform 1 0 1636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1524952243
transform 1 0 1644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1524952243
transform 1 0 1548 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_2756
timestamp 1524952243
transform 1 0 1556 0 1 115
box -3 -3 3 3
use NAND2X1  NAND2X1_50
timestamp 1524952243
transform 1 0 1528 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_2732
timestamp 1524952243
transform 1 0 1660 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1524952243
transform 1 0 1708 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_2377
timestamp 1524952243
transform 1 0 1692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1524952243
transform 1 0 1684 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2757
timestamp 1524952243
transform 1 0 1644 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1524952243
transform 1 0 1668 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1524952243
transform 1 0 1612 0 1 105
box -3 -3 3 3
use XNOR2X1  XNOR2X1_72
timestamp 1524952243
transform -1 0 1608 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2787
timestamp 1524952243
transform 1 0 1636 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_78
timestamp 1524952243
transform 1 0 1608 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_2733
timestamp 1524952243
transform 1 0 1692 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1524952243
transform 1 0 1748 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2378
timestamp 1524952243
transform 1 0 1732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1524952243
transform 1 0 1708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1524952243
transform 1 0 1692 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_2777
timestamp 1524952243
transform 1 0 1684 0 1 105
box -3 -3 3 3
use M2_M1  M2_M1_2457
timestamp 1524952243
transform 1 0 1692 0 1 105
box -2 -2 2 2
use AND2X2  AND2X2_31
timestamp 1524952243
transform -1 0 1696 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_2734
timestamp 1524952243
transform 1 0 1724 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2439
timestamp 1524952243
transform 1 0 1732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1524952243
transform 1 0 1724 0 1 115
box -2 -2 2 2
use NAND3X1  NAND3X1_35
timestamp 1524952243
transform 1 0 1696 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_2684
timestamp 1524952243
transform 1 0 1796 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1524952243
transform 1 0 1828 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1524952243
transform 1 0 1852 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1524952243
transform 1 0 1876 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1524952243
transform 1 0 1780 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1524952243
transform 1 0 1796 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1524952243
transform 1 0 1836 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_2379
timestamp 1524952243
transform 1 0 1780 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1524952243
transform 1 0 1796 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1524952243
transform 1 0 1812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1524952243
transform 1 0 1820 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_2697
timestamp 1524952243
transform 1 0 1884 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1524952243
transform 1 0 1860 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_2440
timestamp 1524952243
transform 1 0 1788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1524952243
transform 1 0 1804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1524952243
transform 1 0 1828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1524952243
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2798
timestamp 1524952243
transform 1 0 1788 0 1 75
box -3 -3 3 3
use XOR2X1  XOR2X1_79
timestamp 1524952243
transform -1 0 1784 0 -1 170
box -8 -3 64 105
use AOI22X1  AOI22X1_93
timestamp 1524952243
transform 1 0 1784 0 -1 170
box -8 -3 46 105
use M2_M1  M2_M1_2383
timestamp 1524952243
transform 1 0 1916 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1524952243
transform 1 0 1892 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1524952243
transform 1 0 1908 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2735
timestamp 1524952243
transform 1 0 1916 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2446
timestamp 1524952243
transform 1 0 1924 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_2736
timestamp 1524952243
transform 1 0 1932 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_2447
timestamp 1524952243
transform 1 0 1940 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1524952243
transform 1 0 1852 0 1 115
box -2 -2 2 2
use OAI21X1  OAI21X1_99
timestamp 1524952243
transform 1 0 1824 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_2759
timestamp 1524952243
transform 1 0 1892 0 1 115
box -3 -3 3 3
use XNOR2X1  XNOR2X1_73
timestamp 1524952243
transform 1 0 1856 0 -1 170
box -8 -3 64 105
use AND2X2  AND2X2_32
timestamp 1524952243
transform 1 0 1912 0 -1 170
box -8 -3 40 105
use top_module_VIA0  top_module_VIA0_37
timestamp 1524952243
transform 1 0 1994 0 1 70
box -10 -3 10 3
use M3_M2  M3_M2_2799
timestamp 1524952243
transform 1 0 972 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1524952243
transform 1 0 1252 0 1 65
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1524952243
transform 1 0 48 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_2801
timestamp 1524952243
transform 1 0 1148 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1524952243
transform 1 0 1284 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1524952243
transform 1 0 964 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1524952243
transform 1 0 1188 0 1 45
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1524952243
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_2805
timestamp 1524952243
transform 1 0 1060 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1524952243
transform 1 0 1220 0 1 35
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1524952243
transform 1 0 1970 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_2807
timestamp 1524952243
transform 1 0 596 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1524952243
transform 1 0 1204 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1524952243
transform 1 0 764 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1524952243
transform 1 0 1084 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1524952243
transform 1 0 1132 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1524952243
transform 1 0 1364 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1524952243
transform 1 0 1396 0 1 15
box -3 -3 3 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1524952243
transform 1 0 1994 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal2 1428 1938 1428 1938 4 in_clka
rlabel metal2 972 1938 972 1938 4 in_clkb
rlabel metal2 604 1938 604 1938 4 in_timer5
rlabel metal2 660 1938 660 1938 4 in_inp
rlabel metal2 588 1938 588 1938 4 in_run
rlabel metal2 876 1938 876 1938 4 in_wai
rlabel metal2 860 1938 860 1938 4 in_reset
rlabel metal3 2 1335 2 1335 4 in_DataIn
rlabel metal3 2 1525 2 1525 4 con_loadData
rlabel metal3 2 1475 2 1475 4 con_readData
rlabel metal2 492 1938 492 1938 4 con_writeData
rlabel metal2 572 1938 572 1938 4 con_writeout
rlabel metal3 2 1035 2 1035 4 con_restart
rlabel metal2 1252 1 1252 1 4 out_MuxData[15]
rlabel metal2 1220 1 1220 1 4 out_MuxData[14]
rlabel metal2 1268 1 1268 1 4 out_MuxData[13]
rlabel metal2 1084 1 1084 1 4 out_MuxData[12]
rlabel metal2 1364 1 1364 1 4 out_MuxData[11]
rlabel metal3 2018 575 2018 575 4 out_MuxData[10]
rlabel metal3 2018 605 2018 605 4 out_MuxData[9]
rlabel metal3 2018 675 2018 675 4 out_MuxData[8]
rlabel metal2 1204 1 1204 1 4 out_MuxData[7]
rlabel metal2 1188 1 1188 1 4 out_MuxData[6]
rlabel metal2 1284 1 1284 1 4 out_MuxData[5]
rlabel metal2 1100 1 1100 1 4 out_MuxData[4]
rlabel metal3 2018 695 2018 695 4 out_MuxData[3]
rlabel metal3 2018 715 2018 715 4 out_MuxData[2]
rlabel metal3 2018 785 2018 785 4 out_MuxData[1]
rlabel metal3 2018 765 2018 765 4 out_MuxData[0]
rlabel metal3 2 365 2 365 4 out_MemBData[15]
rlabel metal3 2 485 2 485 4 out_MemBData[14]
rlabel metal3 2 755 2 755 4 out_MemBData[13]
rlabel metal3 2 855 2 855 4 out_MemBData[12]
rlabel metal3 2 385 2 385 4 out_MemBData[11]
rlabel metal3 2 685 2 685 4 out_MemBData[10]
rlabel metal3 2 875 2 875 4 out_MemBData[9]
rlabel metal3 2 955 2 955 4 out_MemBData[8]
rlabel metal3 2 1175 2 1175 4 out_MemBData[7]
rlabel metal3 2 1055 2 1055 4 out_MemBData[6]
rlabel metal2 844 1938 844 1938 4 out_MemBData[5]
rlabel metal3 2 1315 2 1315 4 out_MemBData[4]
rlabel metal2 956 1938 956 1938 4 out_MemBData[3]
rlabel metal2 940 1938 940 1938 4 out_MemBData[2]
rlabel metal2 924 1938 924 1938 4 out_MemBData[1]
rlabel metal2 908 1938 908 1938 4 out_MemBData[0]
rlabel metal3 2 1815 2 1815 4 out_lose
rlabel metal3 2 1735 2 1735 4 out_win
rlabel metal2 892 1938 892 1938 4 out_state[2]
rlabel metal2 524 1938 524 1938 4 out_state[1]
rlabel metal2 828 1938 828 1938 4 out_state[0]
rlabel metal3 2 1255 2 1255 4 con_count[3]
rlabel metal3 2 1155 2 1155 4 con_count[2]
rlabel metal3 2 1295 2 1295 4 con_count[1]
rlabel metal3 2 1225 2 1225 4 con_count[0]
rlabel metal2 1396 1938 1396 1938 4 con_countWriteout[8]
rlabel metal2 1300 1938 1300 1938 4 con_countWriteout[7]
rlabel metal2 1276 1938 1276 1938 4 con_countWriteout[6]
rlabel metal2 1444 1938 1444 1938 4 con_countWriteout[5]
rlabel metal2 1508 1938 1508 1938 4 con_countWriteout[4]
rlabel metal2 1692 1938 1692 1938 4 con_countWriteout[3]
rlabel metal2 1780 1938 1780 1938 4 con_countWriteout[2]
rlabel metal3 2018 1605 2018 1605 4 con_countWriteout[1]
rlabel metal3 2018 1515 2018 1515 4 con_countWriteout[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>
