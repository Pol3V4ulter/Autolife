magic
tech scmos
timestamp 1524952243
<< m2contact >>
rect -2 -2 2 2
<< end >>
