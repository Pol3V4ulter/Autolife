* SPICE3 file created from top_module.ext - technology: scmos

.option scale=0.3u

M1000 NAND3X1_34/B OAI21X1_91/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=292262 ps=120220
M1001 vdd INVX2_135/Y NAND3X1_34/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 NAND2X1_43/a_9_6# OAI21X1_91/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=151038 ps=69566
M1003 NAND3X1_34/B INVX2_135/Y NAND2X1_43/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 OAI21X1_92/a_9_54# OAI21X1_91/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1005 XNOR2X1_60/A INVX2_135/Y OAI21X1_92/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1006 vdd NAND3X1_34/B XNOR2X1_60/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 gnd OAI21X1_91/A OAI21X1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1008 OAI21X1_92/a_2_6# INVX2_135/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 XNOR2X1_60/A NAND3X1_34/B OAI21X1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 vdd XNOR2X1_60/A XNOR2X1_60/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1011 XNOR2X1_60/a_18_54# XNOR2X1_60/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1012 AOI22X1_99/B XNOR2X1_60/a_2_6# XNOR2X1_60/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1013 XNOR2X1_60/a_35_54# XNOR2X1_60/A AOI22X1_99/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1014 vdd AND2X2_41/Y XNOR2X1_60/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 XNOR2X1_60/a_12_41# AND2X2_41/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1016 gnd XNOR2X1_60/A XNOR2X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1017 XNOR2X1_60/a_18_6# XNOR2X1_60/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1018 AOI22X1_99/B XNOR2X1_60/A XNOR2X1_60/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1019 XNOR2X1_60/a_35_6# XNOR2X1_60/a_2_6# AOI22X1_99/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1020 gnd AND2X2_41/Y XNOR2X1_60/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 XNOR2X1_60/a_12_41# AND2X2_41/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1022 NAND3X1_34/Y AND2X2_41/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1023 vdd NAND3X1_34/B NAND3X1_34/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 NAND3X1_34/Y XOR2X1_91/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 NAND3X1_34/a_9_6# AND2X2_41/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1026 NAND3X1_34/a_14_6# NAND3X1_34/B NAND3X1_34/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1027 NAND3X1_34/Y XOR2X1_91/A NAND3X1_34/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1028 vdd XOR2X1_91/A XOR2X1_91/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1029 XOR2X1_91/a_18_54# XOR2X1_91/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1030 XOR2X1_91/Y XOR2X1_91/A XOR2X1_91/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1031 XOR2X1_91/a_35_54# XOR2X1_91/a_2_6# XOR2X1_91/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1032 vdd AND2X2_41/A XOR2X1_91/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1033 XOR2X1_91/a_13_43# AND2X2_41/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1034 gnd XOR2X1_91/A XOR2X1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1035 XOR2X1_91/a_18_6# XOR2X1_91/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1036 XOR2X1_91/Y XOR2X1_91/a_2_6# XOR2X1_91/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1037 XOR2X1_91/a_35_6# XOR2X1_91/A XOR2X1_91/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1038 gnd AND2X2_41/A XOR2X1_91/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 XOR2X1_91/a_13_43# AND2X2_41/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1040 vdd OAI21X1_90/Y XNOR2X1_59/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1041 XNOR2X1_59/a_18_54# XNOR2X1_59/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1042 AOI22X1_99/D XNOR2X1_59/a_2_6# XNOR2X1_59/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1043 XNOR2X1_59/a_35_54# OAI21X1_90/Y AOI22X1_99/D vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1044 vdd AND2X2_40/Y XNOR2X1_59/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 XNOR2X1_59/a_12_41# AND2X2_40/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1046 gnd OAI21X1_90/Y XNOR2X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1047 XNOR2X1_59/a_18_6# XNOR2X1_59/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1048 AOI22X1_99/D OAI21X1_90/Y XNOR2X1_59/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1049 XNOR2X1_59/a_35_6# XNOR2X1_59/a_2_6# AOI22X1_99/D Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1050 gnd AND2X2_40/Y XNOR2X1_59/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 XNOR2X1_59/a_12_41# AND2X2_40/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1052 vdd XOR2X1_90/A XOR2X1_90/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1053 XOR2X1_90/a_18_54# XOR2X1_90/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1054 XOR2X1_90/Y XOR2X1_90/A XOR2X1_90/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1055 XOR2X1_90/a_35_54# XOR2X1_90/a_2_6# XOR2X1_90/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1056 vdd AND2X2_40/A XOR2X1_90/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 XOR2X1_90/a_13_43# AND2X2_40/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1058 gnd XOR2X1_90/A XOR2X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1059 XOR2X1_90/a_18_6# XOR2X1_90/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1060 XOR2X1_90/Y XOR2X1_90/a_2_6# XOR2X1_90/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1061 XOR2X1_90/a_35_6# XOR2X1_90/A XOR2X1_90/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1062 gnd AND2X2_40/A XOR2X1_90/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 XOR2X1_90/a_13_43# AND2X2_40/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1064 vdd NOR2X1_46/B AOI22X1_99/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1065 AOI22X1_99/a_2_54# AOI22X1_99/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 AOI22X1_99/Y AOI22X1_99/D AOI22X1_99/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1067 AOI22X1_99/a_2_54# NOR2X1_48/B AOI22X1_99/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 AOI22X1_99/a_11_6# NOR2X1_46/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1069 AOI22X1_99/Y AOI22X1_99/B AOI22X1_99/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1070 AOI22X1_99/a_28_6# AOI22X1_99/D AOI22X1_99/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1071 gnd NOR2X1_48/B AOI22X1_99/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 vdd XOR2X1_90/Y AOI22X1_98/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1073 AOI22X1_98/a_2_54# NOR2X1_48/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 AND2X2_38/B NOR2X1_46/B AOI22X1_98/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1075 AOI22X1_98/a_2_54# XOR2X1_91/Y AND2X2_38/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 AOI22X1_98/a_11_6# XOR2X1_90/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1077 AND2X2_38/B NOR2X1_48/B AOI22X1_98/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1078 AOI22X1_98/a_28_6# NOR2X1_46/B AND2X2_38/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1079 gnd XOR2X1_91/Y AOI22X1_98/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 vdd XOR2X1_87/A XOR2X1_87/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1081 XOR2X1_87/a_18_54# XOR2X1_87/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1082 XOR2X1_87/Y XOR2X1_87/A XOR2X1_87/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1083 XOR2X1_87/a_35_54# XOR2X1_87/a_2_6# XOR2X1_87/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1084 vdd XOR2X1_87/B XOR2X1_87/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 XOR2X1_87/a_13_43# XOR2X1_87/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1086 gnd XOR2X1_87/A XOR2X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1087 XOR2X1_87/a_18_6# XOR2X1_87/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1088 XOR2X1_87/Y XOR2X1_87/a_2_6# XOR2X1_87/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1089 XOR2X1_87/a_35_6# XOR2X1_87/A XOR2X1_87/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1090 gnd XOR2X1_87/B XOR2X1_87/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 XOR2X1_87/a_13_43# XOR2X1_87/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1092 AND2X2_38/a_2_6# AND2X2_38/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1093 vdd AND2X2_38/B AND2X2_38/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 AND2X2_38/Y AND2X2_38/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1095 AND2X2_38/a_9_6# AND2X2_38/A AND2X2_38/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1096 gnd AND2X2_38/B AND2X2_38/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 AND2X2_38/Y AND2X2_38/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1098 vdd XOR2X1_86/Y AOI22X1_97/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1099 AOI22X1_97/a_2_54# NOR2X1_47/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 AND2X2_38/A NOR2X1_49/B AOI22X1_97/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1101 AOI22X1_97/a_2_54# XOR2X1_87/Y AND2X2_38/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 AOI22X1_97/a_11_6# XOR2X1_86/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1103 AND2X2_38/A NOR2X1_47/B AOI22X1_97/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1104 AOI22X1_97/a_28_6# NOR2X1_49/B AND2X2_38/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1105 gnd XOR2X1_87/Y AOI22X1_97/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 vdd AND2X2_36/B XOR2X1_86/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1107 XOR2X1_86/a_18_54# XOR2X1_86/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1108 XOR2X1_86/Y AND2X2_36/B XOR2X1_86/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1109 XOR2X1_86/a_35_54# XOR2X1_86/a_2_6# XOR2X1_86/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1110 vdd AND2X2_36/A XOR2X1_86/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 XOR2X1_86/a_13_43# AND2X2_36/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1112 gnd AND2X2_36/B XOR2X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1113 XOR2X1_86/a_18_6# XOR2X1_86/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1114 XOR2X1_86/Y XOR2X1_86/a_2_6# XOR2X1_86/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1115 XOR2X1_86/a_35_6# AND2X2_36/B XOR2X1_86/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1116 gnd AND2X2_36/A XOR2X1_86/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 XOR2X1_86/a_13_43# AND2X2_36/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1118 AND2X2_36/a_2_6# AND2X2_36/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1119 vdd AND2X2_36/B AND2X2_36/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 AND2X2_36/Y AND2X2_36/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1121 AND2X2_36/a_9_6# AND2X2_36/A AND2X2_36/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1122 gnd AND2X2_36/B AND2X2_36/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 AND2X2_36/Y AND2X2_36/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1124 vdd OAI21X1_88/Y XNOR2X1_57/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1125 XNOR2X1_57/a_18_54# XNOR2X1_57/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1126 XNOR2X1_57/Y XNOR2X1_57/a_2_6# XNOR2X1_57/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1127 XNOR2X1_57/a_35_54# OAI21X1_88/Y XNOR2X1_57/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1128 vdd AND2X2_36/Y XNOR2X1_57/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 XNOR2X1_57/a_12_41# AND2X2_36/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1130 gnd OAI21X1_88/Y XNOR2X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1131 XNOR2X1_57/a_18_6# XNOR2X1_57/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1132 XNOR2X1_57/Y OAI21X1_88/Y XNOR2X1_57/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1133 XNOR2X1_57/a_35_6# XNOR2X1_57/a_2_6# XNOR2X1_57/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1134 gnd AND2X2_36/Y XNOR2X1_57/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 XNOR2X1_57/a_12_41# AND2X2_36/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1136 OAI21X1_88/a_9_54# OAI21X1_87/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1137 OAI21X1_88/Y INVX2_123/Y OAI21X1_88/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1138 vdd NAND2X1_42/Y OAI21X1_88/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 gnd OAI21X1_87/A OAI21X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1140 OAI21X1_88/a_2_6# INVX2_123/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 OAI21X1_88/Y NAND2X1_42/Y OAI21X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1142 NAND2X1_42/Y OAI21X1_87/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1143 vdd INVX2_123/Y NAND2X1_42/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 NAND2X1_42/a_9_6# OAI21X1_87/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1145 NAND2X1_42/Y INVX2_123/Y NAND2X1_42/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1146 INVX2_134/Y INVX2_134/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1147 INVX2_134/Y INVX2_134/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1148 vdd INVX2_61/Y DFFPOSX1_100/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1149 DFFPOSX1_100/a_17_74# OAI22X1_19/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1150 DFFPOSX1_100/a_22_6# INVX2_61/Y DFFPOSX1_100/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1151 DFFPOSX1_100/a_31_74# DFFPOSX1_100/a_2_6# DFFPOSX1_100/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1152 vdd DFFPOSX1_100/a_34_4# DFFPOSX1_100/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 DFFPOSX1_100/a_34_4# DFFPOSX1_100/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1154 DFFPOSX1_100/a_61_74# DFFPOSX1_100/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1155 DFFPOSX1_100/a_66_6# DFFPOSX1_100/a_2_6# DFFPOSX1_100/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1156 DFFPOSX1_100/a_76_84# INVX2_61/Y DFFPOSX1_100/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1157 vdd INVX2_134/A DFFPOSX1_100/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 gnd INVX2_61/Y DFFPOSX1_100/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1159 INVX2_134/A DFFPOSX1_100/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1160 DFFPOSX1_100/a_17_6# OAI22X1_19/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1161 DFFPOSX1_100/a_22_6# DFFPOSX1_100/a_2_6# DFFPOSX1_100/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 DFFPOSX1_100/a_31_6# INVX2_61/Y DFFPOSX1_100/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1163 gnd DFFPOSX1_100/a_34_4# DFFPOSX1_100/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 DFFPOSX1_100/a_34_4# DFFPOSX1_100/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1165 DFFPOSX1_100/a_61_6# DFFPOSX1_100/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1166 DFFPOSX1_100/a_66_6# INVX2_61/Y DFFPOSX1_100/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1167 DFFPOSX1_100/a_76_6# DFFPOSX1_100/a_2_6# DFFPOSX1_100/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1168 gnd INVX2_134/A DFFPOSX1_100/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 INVX2_134/A DFFPOSX1_100/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1170 vdd INVX2_61/Y DFFPOSX1_99/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1171 DFFPOSX1_99/a_17_74# OAI22X1_21/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1172 DFFPOSX1_99/a_22_6# INVX2_61/Y DFFPOSX1_99/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1173 DFFPOSX1_99/a_31_74# DFFPOSX1_99/a_2_6# DFFPOSX1_99/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1174 vdd DFFPOSX1_99/a_34_4# DFFPOSX1_99/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 DFFPOSX1_99/a_34_4# DFFPOSX1_99/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1176 DFFPOSX1_99/a_61_74# DFFPOSX1_99/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1177 DFFPOSX1_99/a_66_6# DFFPOSX1_99/a_2_6# DFFPOSX1_99/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1178 DFFPOSX1_99/a_76_84# INVX2_61/Y DFFPOSX1_99/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1179 vdd INVX2_133/A DFFPOSX1_99/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 gnd INVX2_61/Y DFFPOSX1_99/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1181 INVX2_133/A DFFPOSX1_99/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1182 DFFPOSX1_99/a_17_6# OAI22X1_21/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1183 DFFPOSX1_99/a_22_6# DFFPOSX1_99/a_2_6# DFFPOSX1_99/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1184 DFFPOSX1_99/a_31_6# INVX2_61/Y DFFPOSX1_99/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1185 gnd DFFPOSX1_99/a_34_4# DFFPOSX1_99/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 DFFPOSX1_99/a_34_4# DFFPOSX1_99/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1187 DFFPOSX1_99/a_61_6# DFFPOSX1_99/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1188 DFFPOSX1_99/a_66_6# INVX2_61/Y DFFPOSX1_99/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1189 DFFPOSX1_99/a_76_6# DFFPOSX1_99/a_2_6# DFFPOSX1_99/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1190 gnd INVX2_133/A DFFPOSX1_99/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 INVX2_133/A DFFPOSX1_99/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1192 OAI22X1_21/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1193 OAI22X1_21/Y INVX2_133/Y OAI22X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1194 OAI22X1_21/a_28_54# INVX2_131/Y OAI22X1_21/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1195 vdd INVX2_62/Y OAI22X1_21/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 gnd BUFX2_4/Y OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1197 OAI22X1_21/a_2_6# INVX2_133/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 OAI22X1_21/Y INVX2_131/Y OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1199 OAI22X1_21/a_2_6# INVX2_62/Y OAI22X1_21/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 OAI22X1_19/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1201 OAI22X1_19/Y INVX2_134/Y OAI22X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1202 OAI22X1_19/a_28_54# INVX2_129/Y OAI22X1_19/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1203 vdd INVX2_62/Y OAI22X1_19/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 gnd BUFX2_4/Y OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1205 OAI22X1_19/a_2_6# INVX2_134/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 OAI22X1_19/Y INVX2_129/Y OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1207 OAI22X1_19/a_2_6# INVX2_62/Y OAI22X1_19/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 INVX2_131/Y out_MemBData[7] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1209 INVX2_131/Y out_MemBData[7] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1210 NOR2X1_49/a_9_54# INVX2_62/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1211 NOR2X1_49/Y NOR2X1_49/B NOR2X1_49/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1212 NOR2X1_49/Y INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1213 gnd NOR2X1_49/B NOR2X1_49/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 OAI21X1_86/a_9_54# NOR2X1_49/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1215 OAI21X1_85/C AND2X2_19/Y OAI21X1_86/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1216 vdd out_MemBData[7] OAI21X1_85/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 gnd NOR2X1_49/Y OAI21X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1218 OAI21X1_86/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 OAI21X1_85/C out_MemBData[7] OAI21X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1220 OAI21X1_85/a_9_54# INVX2_130/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1221 OAI21X1_85/Y OR2X2_0/Y OAI21X1_85/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1222 vdd OAI21X1_85/C OAI21X1_85/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 gnd INVX2_130/A OAI21X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1224 OAI21X1_85/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 OAI21X1_85/Y OAI21X1_85/C OAI21X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1226 INVX2_129/Y out_MemBData[6] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1227 INVX2_129/Y out_MemBData[6] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1228 NOR2X1_47/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1229 NOR2X1_47/Y NOR2X1_47/B NOR2X1_47/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1230 NOR2X1_47/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1231 gnd NOR2X1_47/B NOR2X1_47/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 OAI21X1_82/a_9_54# NOR2X1_47/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1233 OAI21X1_80/C AND2X2_19/Y OAI21X1_82/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1234 vdd out_MemBData[6] OAI21X1_80/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 gnd NOR2X1_47/Y OAI21X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1236 OAI21X1_82/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 OAI21X1_80/C out_MemBData[6] OAI21X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1238 OAI21X1_80/a_9_54# INVX2_128/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1239 OAI21X1_80/Y OR2X2_0/Y OAI21X1_80/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1240 vdd OAI21X1_80/C OAI21X1_80/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 gnd INVX2_128/A OAI21X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1242 OAI21X1_80/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 OAI21X1_80/Y OAI21X1_80/C OAI21X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1244 vdd BUFX2_11/Y DFFPOSX1_95/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1245 DFFPOSX1_95/a_17_74# OAI21X1_80/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1246 DFFPOSX1_95/a_22_6# BUFX2_11/Y DFFPOSX1_95/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1247 DFFPOSX1_95/a_31_74# DFFPOSX1_95/a_2_6# DFFPOSX1_95/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1248 vdd DFFPOSX1_95/a_34_4# DFFPOSX1_95/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 DFFPOSX1_95/a_34_4# DFFPOSX1_95/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1250 DFFPOSX1_95/a_61_74# DFFPOSX1_95/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1251 DFFPOSX1_95/a_66_6# DFFPOSX1_95/a_2_6# DFFPOSX1_95/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1252 DFFPOSX1_95/a_76_84# BUFX2_11/Y DFFPOSX1_95/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1253 vdd out_MemBData[6] DFFPOSX1_95/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 gnd BUFX2_11/Y DFFPOSX1_95/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1255 out_MemBData[6] DFFPOSX1_95/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1256 DFFPOSX1_95/a_17_6# OAI21X1_80/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1257 DFFPOSX1_95/a_22_6# DFFPOSX1_95/a_2_6# DFFPOSX1_95/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1258 DFFPOSX1_95/a_31_6# BUFX2_11/Y DFFPOSX1_95/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1259 gnd DFFPOSX1_95/a_34_4# DFFPOSX1_95/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 DFFPOSX1_95/a_34_4# DFFPOSX1_95/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1261 DFFPOSX1_95/a_61_6# DFFPOSX1_95/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1262 DFFPOSX1_95/a_66_6# BUFX2_11/Y DFFPOSX1_95/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1263 DFFPOSX1_95/a_76_6# DFFPOSX1_95/a_2_6# DFFPOSX1_95/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1264 gnd out_MemBData[6] DFFPOSX1_95/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 out_MemBData[6] DFFPOSX1_95/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1266 vdd INVX2_43/Y DFFPOSX1_94/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1267 DFFPOSX1_94/a_17_74# INVX2_127/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1268 DFFPOSX1_94/a_22_6# INVX2_43/Y DFFPOSX1_94/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1269 DFFPOSX1_94/a_31_74# DFFPOSX1_94/a_2_6# DFFPOSX1_94/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1270 vdd DFFPOSX1_94/a_34_4# DFFPOSX1_94/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 DFFPOSX1_94/a_34_4# DFFPOSX1_94/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1272 DFFPOSX1_94/a_61_74# DFFPOSX1_94/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1273 DFFPOSX1_94/a_66_6# DFFPOSX1_94/a_2_6# DFFPOSX1_94/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1274 DFFPOSX1_94/a_76_84# INVX2_43/Y DFFPOSX1_94/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1275 vdd con_count[3] DFFPOSX1_94/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 gnd INVX2_43/Y DFFPOSX1_94/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1277 con_count[3] DFFPOSX1_94/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1278 DFFPOSX1_94/a_17_6# INVX2_127/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1279 DFFPOSX1_94/a_22_6# DFFPOSX1_94/a_2_6# DFFPOSX1_94/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1280 DFFPOSX1_94/a_31_6# INVX2_43/Y DFFPOSX1_94/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1281 gnd DFFPOSX1_94/a_34_4# DFFPOSX1_94/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 DFFPOSX1_94/a_34_4# DFFPOSX1_94/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1283 DFFPOSX1_94/a_61_6# DFFPOSX1_94/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1284 DFFPOSX1_94/a_66_6# INVX2_43/Y DFFPOSX1_94/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1285 DFFPOSX1_94/a_76_6# DFFPOSX1_94/a_2_6# DFFPOSX1_94/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1286 gnd con_count[3] DFFPOSX1_94/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 con_count[3] DFFPOSX1_94/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1288 INVX2_127/Y INVX2_127/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1289 INVX2_127/Y INVX2_127/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1290 vdd BUFX2_9/Y DFFPOSX1_92/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1291 DFFPOSX1_92/a_17_74# AND2X2_34/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1292 DFFPOSX1_92/a_22_6# BUFX2_9/Y DFFPOSX1_92/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1293 DFFPOSX1_92/a_31_74# DFFPOSX1_92/a_2_6# DFFPOSX1_92/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1294 vdd DFFPOSX1_92/a_34_4# DFFPOSX1_92/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 DFFPOSX1_92/a_34_4# DFFPOSX1_92/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1296 DFFPOSX1_92/a_61_74# DFFPOSX1_92/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1297 DFFPOSX1_92/a_66_6# DFFPOSX1_92/a_2_6# DFFPOSX1_92/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1298 DFFPOSX1_92/a_76_84# BUFX2_9/Y DFFPOSX1_92/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1299 vdd AOI22X1_93/C DFFPOSX1_92/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 gnd BUFX2_9/Y DFFPOSX1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1301 AOI22X1_93/C DFFPOSX1_92/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1302 DFFPOSX1_92/a_17_6# AND2X2_34/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1303 DFFPOSX1_92/a_22_6# DFFPOSX1_92/a_2_6# DFFPOSX1_92/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1304 DFFPOSX1_92/a_31_6# BUFX2_9/Y DFFPOSX1_92/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1305 gnd DFFPOSX1_92/a_34_4# DFFPOSX1_92/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1306 DFFPOSX1_92/a_34_4# DFFPOSX1_92/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1307 DFFPOSX1_92/a_61_6# DFFPOSX1_92/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1308 DFFPOSX1_92/a_66_6# BUFX2_9/Y DFFPOSX1_92/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1309 DFFPOSX1_92/a_76_6# DFFPOSX1_92/a_2_6# DFFPOSX1_92/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1310 gnd AOI22X1_93/C DFFPOSX1_92/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 AOI22X1_93/C DFFPOSX1_92/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1312 INVX2_125/Y INVX2_125/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1313 INVX2_125/Y INVX2_125/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1314 vdd INVX2_43/Y DFFPOSX1_91/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1315 DFFPOSX1_91/a_17_74# INVX2_125/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1316 DFFPOSX1_91/a_22_6# INVX2_43/Y DFFPOSX1_91/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1317 DFFPOSX1_91/a_31_74# DFFPOSX1_91/a_2_6# DFFPOSX1_91/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1318 vdd DFFPOSX1_91/a_34_4# DFFPOSX1_91/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 DFFPOSX1_91/a_34_4# DFFPOSX1_91/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1320 DFFPOSX1_91/a_61_74# DFFPOSX1_91/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1321 DFFPOSX1_91/a_66_6# DFFPOSX1_91/a_2_6# DFFPOSX1_91/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1322 DFFPOSX1_91/a_76_84# INVX2_43/Y DFFPOSX1_91/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1323 vdd con_count[4] DFFPOSX1_91/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1324 gnd INVX2_43/Y DFFPOSX1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1325 con_count[4] DFFPOSX1_91/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1326 DFFPOSX1_91/a_17_6# INVX2_125/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1327 DFFPOSX1_91/a_22_6# DFFPOSX1_91/a_2_6# DFFPOSX1_91/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1328 DFFPOSX1_91/a_31_6# INVX2_43/Y DFFPOSX1_91/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1329 gnd DFFPOSX1_91/a_34_4# DFFPOSX1_91/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 DFFPOSX1_91/a_34_4# DFFPOSX1_91/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1331 DFFPOSX1_91/a_61_6# DFFPOSX1_91/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1332 DFFPOSX1_91/a_66_6# INVX2_43/Y DFFPOSX1_91/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1333 DFFPOSX1_91/a_76_6# DFFPOSX1_91/a_2_6# DFFPOSX1_91/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1334 gnd con_count[4] DFFPOSX1_91/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 con_count[4] DFFPOSX1_91/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1336 INVX2_135/Y INVX2_135/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1337 INVX2_135/Y INVX2_135/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1338 OAI21X1_91/a_9_54# OAI21X1_91/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1339 XOR2X1_89/A INVX2_135/Y OAI21X1_91/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1340 vdd NAND3X1_34/Y XOR2X1_89/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1341 gnd OAI21X1_91/A OAI21X1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1342 OAI21X1_91/a_2_6# INVX2_135/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 XOR2X1_89/A NAND3X1_34/Y OAI21X1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1344 vdd XOR2X1_89/A XOR2X1_89/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1345 XOR2X1_89/a_18_54# XOR2X1_89/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1346 XOR2X1_89/Y XOR2X1_89/A XOR2X1_89/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1347 XOR2X1_89/a_35_54# XOR2X1_89/a_2_6# XOR2X1_89/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1348 vdd XOR2X1_89/B XOR2X1_89/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 XOR2X1_89/a_13_43# XOR2X1_89/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1350 gnd XOR2X1_89/A XOR2X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1351 XOR2X1_89/a_18_6# XOR2X1_89/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1352 XOR2X1_89/Y XOR2X1_89/a_2_6# XOR2X1_89/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1353 XOR2X1_89/a_35_6# XOR2X1_89/A XOR2X1_89/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1354 gnd XOR2X1_89/B XOR2X1_89/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 XOR2X1_89/a_13_43# XOR2X1_89/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1356 AND2X2_41/a_2_6# AND2X2_41/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1357 vdd XOR2X1_91/A AND2X2_41/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 AND2X2_41/Y AND2X2_41/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1359 AND2X2_41/a_9_6# AND2X2_41/A AND2X2_41/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1360 gnd XOR2X1_91/A AND2X2_41/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1361 AND2X2_41/Y AND2X2_41/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1362 OAI21X1_90/a_9_54# OAI21X1_89/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1363 OAI21X1_90/Y OAI21X1_89/B OAI21X1_90/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1364 vdd OAI21X1_90/C OAI21X1_90/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 gnd OAI21X1_89/A OAI21X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1366 OAI21X1_90/a_2_6# OAI21X1_89/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 OAI21X1_90/Y OAI21X1_90/C OAI21X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1368 AND2X2_40/a_2_6# AND2X2_40/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1369 vdd XOR2X1_90/A AND2X2_40/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1370 AND2X2_40/Y AND2X2_40/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1371 AND2X2_40/a_9_6# AND2X2_40/A AND2X2_40/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1372 gnd XOR2X1_90/A AND2X2_40/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1373 AND2X2_40/Y AND2X2_40/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1374 OAI21X1_89/a_9_54# OAI21X1_89/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1375 XOR2X1_88/A OAI21X1_89/B OAI21X1_89/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1376 vdd OAI21X1_89/C XOR2X1_88/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 gnd OAI21X1_89/A OAI21X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1378 OAI21X1_89/a_2_6# OAI21X1_89/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 XOR2X1_88/A OAI21X1_89/C OAI21X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1380 vdd XOR2X1_88/A XOR2X1_88/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1381 XOR2X1_88/a_18_54# XOR2X1_88/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1382 XOR2X1_88/Y XOR2X1_88/A XOR2X1_88/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1383 XOR2X1_88/a_35_54# XOR2X1_88/a_2_6# XOR2X1_88/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1384 vdd XOR2X1_88/B XOR2X1_88/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1385 XOR2X1_88/a_13_43# XOR2X1_88/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1386 gnd XOR2X1_88/A XOR2X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1387 XOR2X1_88/a_18_6# XOR2X1_88/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1388 XOR2X1_88/Y XOR2X1_88/a_2_6# XOR2X1_88/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1389 XOR2X1_88/a_35_6# XOR2X1_88/A XOR2X1_88/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1390 gnd XOR2X1_88/B XOR2X1_88/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 XOR2X1_88/a_13_43# XOR2X1_88/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1392 AND2X2_39/a_2_6# AND2X2_39/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1393 vdd AND2X2_39/B AND2X2_39/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 AND2X2_39/Y AND2X2_39/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1395 AND2X2_39/a_9_6# AND2X2_39/A AND2X2_39/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1396 gnd AND2X2_39/B AND2X2_39/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1397 AND2X2_39/Y AND2X2_39/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1398 AND2X2_37/a_2_6# XOR2X1_87/B vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1399 vdd XOR2X1_87/A AND2X2_37/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 AND2X2_37/Y AND2X2_37/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1401 AND2X2_37/a_9_6# XOR2X1_87/B AND2X2_37/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1402 gnd XOR2X1_87/A AND2X2_37/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 AND2X2_37/Y AND2X2_37/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1404 vdd XNOR2X1_58/A XNOR2X1_58/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1405 XNOR2X1_58/a_18_54# XNOR2X1_58/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1406 AOI22X1_96/B XNOR2X1_58/a_2_6# XNOR2X1_58/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1407 XNOR2X1_58/a_35_54# XNOR2X1_58/A AOI22X1_96/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1408 vdd AND2X2_37/Y XNOR2X1_58/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 XNOR2X1_58/a_12_41# AND2X2_37/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1410 gnd XNOR2X1_58/A XNOR2X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1411 XNOR2X1_58/a_18_6# XNOR2X1_58/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1412 AOI22X1_96/B XNOR2X1_58/A XNOR2X1_58/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1413 XNOR2X1_58/a_35_6# XNOR2X1_58/a_2_6# AOI22X1_96/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1414 gnd AND2X2_37/Y XNOR2X1_58/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 XNOR2X1_58/a_12_41# AND2X2_37/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1416 vdd NOR2X1_49/B AOI22X1_96/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1417 AOI22X1_96/a_2_54# AOI22X1_96/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1418 AOI22X1_96/Y XNOR2X1_57/Y AOI22X1_96/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1419 AOI22X1_96/a_2_54# NOR2X1_47/B AOI22X1_96/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1420 AOI22X1_96/a_11_6# NOR2X1_49/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1421 AOI22X1_96/Y AOI22X1_96/B AOI22X1_96/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1422 AOI22X1_96/a_28_6# XNOR2X1_57/Y AOI22X1_96/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1423 gnd NOR2X1_47/B AOI22X1_96/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 vdd XOR2X1_85/Y AOI22X1_95/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1425 AOI22X1_95/a_2_54# NOR2X1_47/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 AND2X2_39/A NOR2X1_49/B AOI22X1_95/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1427 AOI22X1_95/a_2_54# XOR2X1_82/Y AND2X2_39/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 AOI22X1_95/a_11_6# XOR2X1_85/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1429 AND2X2_39/A NOR2X1_47/B AOI22X1_95/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1430 AOI22X1_95/a_28_6# NOR2X1_49/B AND2X2_39/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1431 gnd XOR2X1_82/Y AOI22X1_95/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 vdd XOR2X1_85/A XOR2X1_85/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1433 XOR2X1_85/a_18_54# XOR2X1_85/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1434 XOR2X1_85/Y XOR2X1_85/A XOR2X1_85/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1435 XOR2X1_85/a_35_54# XOR2X1_85/a_2_6# XOR2X1_85/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1436 vdd XOR2X1_85/B XOR2X1_85/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1437 XOR2X1_85/a_13_43# XOR2X1_85/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1438 gnd XOR2X1_85/A XOR2X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1439 XOR2X1_85/a_18_6# XOR2X1_85/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1440 XOR2X1_85/Y XOR2X1_85/a_2_6# XOR2X1_85/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1441 XOR2X1_85/a_35_6# XOR2X1_85/A XOR2X1_85/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1442 gnd XOR2X1_85/B XOR2X1_85/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1443 XOR2X1_85/a_13_43# XOR2X1_85/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1444 OAI21X1_87/C AND2X2_36/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1445 vdd NAND2X1_42/Y OAI21X1_87/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 OAI21X1_87/C AND2X2_36/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 NAND3X1_33/a_9_6# AND2X2_36/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1448 NAND3X1_33/a_14_6# NAND2X1_42/Y NAND3X1_33/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1449 OAI21X1_87/C AND2X2_36/B NAND3X1_33/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1450 OAI21X1_87/a_9_54# OAI21X1_87/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1451 XOR2X1_85/A INVX2_123/Y OAI21X1_87/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1452 vdd OAI21X1_87/C XOR2X1_85/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 gnd OAI21X1_87/A OAI21X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1454 OAI21X1_87/a_2_6# INVX2_123/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 XOR2X1_85/A OAI21X1_87/C OAI21X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1456 vdd BUFX2_10/Y DFFPOSX1_98/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1457 DFFPOSX1_98/a_17_74# OAI22X1_17/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1458 DFFPOSX1_98/a_22_6# BUFX2_10/Y DFFPOSX1_98/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1459 DFFPOSX1_98/a_31_74# DFFPOSX1_98/a_2_6# DFFPOSX1_98/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1460 vdd DFFPOSX1_98/a_34_4# DFFPOSX1_98/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 DFFPOSX1_98/a_34_4# DFFPOSX1_98/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1462 DFFPOSX1_98/a_61_74# DFFPOSX1_98/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1463 DFFPOSX1_98/a_66_6# DFFPOSX1_98/a_2_6# DFFPOSX1_98/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1464 DFFPOSX1_98/a_76_84# BUFX2_10/Y DFFPOSX1_98/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1465 vdd out_MuxData[11] DFFPOSX1_98/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 gnd BUFX2_10/Y DFFPOSX1_98/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1467 out_MuxData[11] DFFPOSX1_98/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1468 DFFPOSX1_98/a_17_6# OAI22X1_17/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1469 DFFPOSX1_98/a_22_6# DFFPOSX1_98/a_2_6# DFFPOSX1_98/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1470 DFFPOSX1_98/a_31_6# BUFX2_10/Y DFFPOSX1_98/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1471 gnd DFFPOSX1_98/a_34_4# DFFPOSX1_98/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 DFFPOSX1_98/a_34_4# DFFPOSX1_98/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1473 DFFPOSX1_98/a_61_6# DFFPOSX1_98/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1474 DFFPOSX1_98/a_66_6# BUFX2_10/Y DFFPOSX1_98/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1475 DFFPOSX1_98/a_76_6# DFFPOSX1_98/a_2_6# DFFPOSX1_98/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1476 gnd out_MuxData[11] DFFPOSX1_98/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 out_MuxData[11] DFFPOSX1_98/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1478 INVX2_133/Y INVX2_133/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1479 INVX2_133/Y INVX2_133/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1480 vdd INVX2_61/Y DFFPOSX1_97/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1481 DFFPOSX1_97/a_17_74# OAI22X1_20/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1482 DFFPOSX1_97/a_22_6# INVX2_61/Y DFFPOSX1_97/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1483 DFFPOSX1_97/a_31_74# DFFPOSX1_97/a_2_6# DFFPOSX1_97/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1484 vdd DFFPOSX1_97/a_34_4# DFFPOSX1_97/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 DFFPOSX1_97/a_34_4# DFFPOSX1_97/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1486 DFFPOSX1_97/a_61_74# DFFPOSX1_97/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1487 DFFPOSX1_97/a_66_6# DFFPOSX1_97/a_2_6# DFFPOSX1_97/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1488 DFFPOSX1_97/a_76_84# INVX2_61/Y DFFPOSX1_97/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1489 vdd INVX2_122/A DFFPOSX1_97/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1490 gnd INVX2_61/Y DFFPOSX1_97/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1491 INVX2_122/A DFFPOSX1_97/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1492 DFFPOSX1_97/a_17_6# OAI22X1_20/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1493 DFFPOSX1_97/a_22_6# DFFPOSX1_97/a_2_6# DFFPOSX1_97/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1494 DFFPOSX1_97/a_31_6# INVX2_61/Y DFFPOSX1_97/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1495 gnd DFFPOSX1_97/a_34_4# DFFPOSX1_97/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 DFFPOSX1_97/a_34_4# DFFPOSX1_97/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1497 DFFPOSX1_97/a_61_6# DFFPOSX1_97/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1498 DFFPOSX1_97/a_66_6# INVX2_61/Y DFFPOSX1_97/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1499 DFFPOSX1_97/a_76_6# DFFPOSX1_97/a_2_6# DFFPOSX1_97/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1500 gnd INVX2_122/A DFFPOSX1_97/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 INVX2_122/A DFFPOSX1_97/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1502 OAI22X1_20/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1503 OAI22X1_20/Y INVX2_122/Y OAI22X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1504 OAI22X1_20/a_28_54# INVX2_132/Y OAI22X1_20/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1505 vdd INVX2_62/Y OAI22X1_20/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 gnd BUFX2_4/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1507 OAI22X1_20/a_2_6# INVX2_122/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1508 OAI22X1_20/Y INVX2_132/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1509 OAI22X1_20/a_2_6# INVX2_62/Y OAI22X1_20/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 INVX2_132/Y out_MemBData[11] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1511 INVX2_132/Y out_MemBData[11] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1512 NOR2X1_49/B INVX2_130/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1513 NOR2X1_49/B INVX2_130/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1514 vdd BUFX2_10/Y DFFPOSX1_96/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1515 DFFPOSX1_96/a_17_74# OAI21X1_85/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1516 DFFPOSX1_96/a_22_6# BUFX2_10/Y DFFPOSX1_96/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1517 DFFPOSX1_96/a_31_74# DFFPOSX1_96/a_2_6# DFFPOSX1_96/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1518 vdd DFFPOSX1_96/a_34_4# DFFPOSX1_96/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1519 DFFPOSX1_96/a_34_4# DFFPOSX1_96/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1520 DFFPOSX1_96/a_61_74# DFFPOSX1_96/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1521 DFFPOSX1_96/a_66_6# DFFPOSX1_96/a_2_6# DFFPOSX1_96/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1522 DFFPOSX1_96/a_76_84# BUFX2_10/Y DFFPOSX1_96/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1523 vdd out_MemBData[7] DFFPOSX1_96/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 gnd BUFX2_10/Y DFFPOSX1_96/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1525 out_MemBData[7] DFFPOSX1_96/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1526 DFFPOSX1_96/a_17_6# OAI21X1_85/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1527 DFFPOSX1_96/a_22_6# DFFPOSX1_96/a_2_6# DFFPOSX1_96/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1528 DFFPOSX1_96/a_31_6# BUFX2_10/Y DFFPOSX1_96/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1529 gnd DFFPOSX1_96/a_34_4# DFFPOSX1_96/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 DFFPOSX1_96/a_34_4# DFFPOSX1_96/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1531 DFFPOSX1_96/a_61_6# DFFPOSX1_96/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1532 DFFPOSX1_96/a_66_6# BUFX2_10/Y DFFPOSX1_96/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1533 DFFPOSX1_96/a_76_6# DFFPOSX1_96/a_2_6# DFFPOSX1_96/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1534 gnd out_MemBData[7] DFFPOSX1_96/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1535 out_MemBData[7] DFFPOSX1_96/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1536 NOR2X1_48/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1537 NOR2X1_48/Y NOR2X1_48/B NOR2X1_48/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1538 NOR2X1_48/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1539 gnd NOR2X1_48/B NOR2X1_48/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1540 OAI21X1_84/a_9_54# NOR2X1_48/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1541 OAI21X1_84/Y AND2X2_19/Y OAI21X1_84/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1542 vdd out_MemBData[4] OAI21X1_84/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1543 gnd NOR2X1_48/Y OAI21X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1544 OAI21X1_84/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 OAI21X1_84/Y out_MemBData[4] OAI21X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1546 OAI21X1_83/a_9_54# INVX2_118/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1547 OAI21X1_83/Y OR2X2_0/Y OAI21X1_83/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1548 vdd OAI21X1_84/Y OAI21X1_83/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 gnd INVX2_118/A OAI21X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1550 OAI21X1_83/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1551 OAI21X1_83/Y OAI21X1_84/Y OAI21X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1552 OAI21X1_81/a_9_54# NOR2X1_46/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1553 OAI21X1_81/Y AND2X2_19/Y OAI21X1_81/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1554 vdd out_MemBData[5] OAI21X1_81/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1555 gnd NOR2X1_46/Y OAI21X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1556 OAI21X1_81/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 OAI21X1_81/Y out_MemBData[5] OAI21X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1558 NOR2X1_47/B INVX2_128/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1559 NOR2X1_47/B INVX2_128/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1560 NOR2X1_46/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1561 NOR2X1_46/Y NOR2X1_46/B NOR2X1_46/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1562 NOR2X1_46/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1563 gnd NOR2X1_46/B NOR2X1_46/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 vdd BUFX2_9/Y DFFPOSX1_93/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1565 DFFPOSX1_93/a_17_74# AND2X2_35/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1566 DFFPOSX1_93/a_22_6# BUFX2_9/Y DFFPOSX1_93/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1567 DFFPOSX1_93/a_31_74# DFFPOSX1_93/a_2_6# DFFPOSX1_93/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1568 vdd DFFPOSX1_93/a_34_4# DFFPOSX1_93/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 DFFPOSX1_93/a_34_4# DFFPOSX1_93/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1570 DFFPOSX1_93/a_61_74# DFFPOSX1_93/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1571 DFFPOSX1_93/a_66_6# DFFPOSX1_93/a_2_6# DFFPOSX1_93/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1572 DFFPOSX1_93/a_76_84# BUFX2_9/Y DFFPOSX1_93/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1573 vdd AOI22X1_94/C DFFPOSX1_93/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1574 gnd BUFX2_9/Y DFFPOSX1_93/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1575 AOI22X1_94/C DFFPOSX1_93/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1576 DFFPOSX1_93/a_17_6# AND2X2_35/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1577 DFFPOSX1_93/a_22_6# DFFPOSX1_93/a_2_6# DFFPOSX1_93/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1578 DFFPOSX1_93/a_31_6# BUFX2_9/Y DFFPOSX1_93/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1579 gnd DFFPOSX1_93/a_34_4# DFFPOSX1_93/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1580 DFFPOSX1_93/a_34_4# DFFPOSX1_93/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1581 DFFPOSX1_93/a_61_6# DFFPOSX1_93/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1582 DFFPOSX1_93/a_66_6# BUFX2_9/Y DFFPOSX1_93/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1583 DFFPOSX1_93/a_76_6# DFFPOSX1_93/a_2_6# DFFPOSX1_93/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1584 gnd AOI22X1_94/C DFFPOSX1_93/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 AOI22X1_94/C DFFPOSX1_93/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1586 vdd con_count[3] AOI22X1_94/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1587 AOI22X1_94/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1588 INVX2_127/A INVX2_126/A AOI22X1_94/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1589 AOI22X1_94/a_2_54# AOI22X1_94/C INVX2_127/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1590 AOI22X1_94/a_11_6# con_count[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1591 INVX2_127/A INVX2_126/Y AOI22X1_94/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1592 AOI22X1_94/a_28_6# INVX2_126/A INVX2_127/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1593 gnd AOI22X1_94/C AOI22X1_94/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1594 AND2X2_35/a_2_6# HAX1_13/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1595 vdd INVX2_72/Y AND2X2_35/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 AND2X2_35/Y AND2X2_35/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1597 AND2X2_35/a_9_6# HAX1_13/YS AND2X2_35/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1598 gnd INVX2_72/Y AND2X2_35/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1599 AND2X2_35/Y AND2X2_35/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1600 vdd con_count[4] AOI22X1_93/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1601 AOI22X1_93/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1602 INVX2_125/A INVX2_126/A AOI22X1_93/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1603 AOI22X1_93/a_2_54# AOI22X1_93/C INVX2_125/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1604 AOI22X1_93/a_11_6# con_count[4] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1605 INVX2_125/A INVX2_126/Y AOI22X1_93/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1606 AOI22X1_93/a_28_6# INVX2_126/A INVX2_125/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1607 gnd AOI22X1_93/C AOI22X1_93/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1608 AND2X2_34/a_2_6# HAX1_12/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1609 vdd INVX2_72/Y AND2X2_34/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1610 AND2X2_34/Y AND2X2_34/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1611 AND2X2_34/a_9_6# HAX1_12/YS AND2X2_34/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M1612 gnd INVX2_72/Y AND2X2_34/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 AND2X2_34/Y AND2X2_34/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1614 INVX2_126/Y INVX2_126/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1615 INVX2_126/Y INVX2_126/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1616 vdd INVX2_43/Y DFFPOSX1_90/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1617 DFFPOSX1_90/a_17_74# INVX2_124/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1618 DFFPOSX1_90/a_22_6# INVX2_43/Y DFFPOSX1_90/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1619 DFFPOSX1_90/a_31_74# DFFPOSX1_90/a_2_6# DFFPOSX1_90/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1620 vdd DFFPOSX1_90/a_34_4# DFFPOSX1_90/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 DFFPOSX1_90/a_34_4# DFFPOSX1_90/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1622 DFFPOSX1_90/a_61_74# DFFPOSX1_90/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1623 DFFPOSX1_90/a_66_6# DFFPOSX1_90/a_2_6# DFFPOSX1_90/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1624 DFFPOSX1_90/a_76_84# INVX2_43/Y DFFPOSX1_90/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1625 vdd con_count[5] DFFPOSX1_90/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1626 gnd INVX2_43/Y DFFPOSX1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1627 con_count[5] DFFPOSX1_90/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1628 DFFPOSX1_90/a_17_6# INVX2_124/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1629 DFFPOSX1_90/a_22_6# DFFPOSX1_90/a_2_6# DFFPOSX1_90/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1630 DFFPOSX1_90/a_31_6# INVX2_43/Y DFFPOSX1_90/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1631 gnd DFFPOSX1_90/a_34_4# DFFPOSX1_90/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1632 DFFPOSX1_90/a_34_4# DFFPOSX1_90/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1633 DFFPOSX1_90/a_61_6# DFFPOSX1_90/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1634 DFFPOSX1_90/a_66_6# INVX2_43/Y DFFPOSX1_90/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1635 DFFPOSX1_90/a_76_6# DFFPOSX1_90/a_2_6# DFFPOSX1_90/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1636 gnd con_count[5] DFFPOSX1_90/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 con_count[5] DFFPOSX1_90/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1638 INVX2_124/Y INVX2_124/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1639 INVX2_124/Y INVX2_124/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1640 vdd NOR2X1_45/A AOI21X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M1641 AOI21X1_8/a_2_54# NOR2X1_45/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1642 INVX2_135/A XOR2X1_89/B AOI21X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1643 AOI21X1_8/a_12_6# NOR2X1_45/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1644 INVX2_135/A NOR2X1_45/B AOI21X1_8/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M1645 gnd XOR2X1_89/B INVX2_135/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1646 NOR2X1_45/a_9_54# NOR2X1_45/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1647 XOR2X1_89/B NOR2X1_45/B NOR2X1_45/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1648 XOR2X1_89/B NOR2X1_45/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1649 gnd NOR2X1_45/B XOR2X1_89/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1650 vdd XOR2X1_81/A XNOR2X1_56/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1651 XNOR2X1_56/a_18_54# XNOR2X1_56/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1652 AND2X2_41/A XNOR2X1_56/a_2_6# XNOR2X1_56/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1653 XNOR2X1_56/a_35_54# XOR2X1_81/A AND2X2_41/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1654 vdd XOR2X1_83/Y XNOR2X1_56/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1655 XNOR2X1_56/a_12_41# XOR2X1_83/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1656 gnd XOR2X1_81/A XNOR2X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1657 XNOR2X1_56/a_18_6# XNOR2X1_56/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1658 AND2X2_41/A XOR2X1_81/A XNOR2X1_56/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1659 XNOR2X1_56/a_35_6# XNOR2X1_56/a_2_6# AND2X2_41/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1660 gnd XOR2X1_83/Y XNOR2X1_56/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 XNOR2X1_56/a_12_41# XOR2X1_83/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1662 OAI21X1_90/C OAI21X1_89/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1663 vdd OAI21X1_89/B OAI21X1_90/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 NAND2X1_41/a_9_6# OAI21X1_89/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1665 OAI21X1_90/C OAI21X1_89/B NAND2X1_41/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1666 OAI21X1_89/C AND2X2_40/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1667 vdd OAI21X1_90/C OAI21X1_89/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1668 OAI21X1_89/C XOR2X1_90/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 NAND3X1_32/a_9_6# AND2X2_40/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1670 NAND3X1_32/a_14_6# OAI21X1_90/C NAND3X1_32/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1671 OAI21X1_89/C XOR2X1_90/A NAND3X1_32/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1672 NOR2X1_44/a_9_54# NOR2X1_44/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1673 XOR2X1_88/B NOR2X1_44/B NOR2X1_44/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1674 XOR2X1_88/B NOR2X1_44/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1675 gnd NOR2X1_44/B XOR2X1_88/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1676 vdd XOR2X1_88/Y AOI22X1_91/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1677 AOI22X1_91/a_2_54# NOR2X1_48/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1678 AND2X2_39/B NOR2X1_46/B AOI22X1_91/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1679 AOI22X1_91/a_2_54# XOR2X1_89/Y AND2X2_39/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 AOI22X1_91/a_11_6# XOR2X1_88/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1681 AND2X2_39/B NOR2X1_48/B AOI22X1_91/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1682 AOI22X1_91/a_28_6# NOR2X1_46/B AND2X2_39/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1683 gnd XOR2X1_89/Y AOI22X1_91/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1684 OAI21X1_78/C XOR2X1_87/B vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1685 vdd OAI21X1_79/C OAI21X1_78/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1686 OAI21X1_78/C XOR2X1_87/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1687 NAND3X1_31/a_9_6# XOR2X1_87/B gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1688 NAND3X1_31/a_14_6# OAI21X1_79/C NAND3X1_31/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M1689 OAI21X1_78/C XOR2X1_87/A NAND3X1_31/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1690 OAI21X1_79/a_9_54# OAI21X1_78/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1691 XNOR2X1_58/A OAI21X1_78/B OAI21X1_79/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1692 vdd OAI21X1_79/C XNOR2X1_58/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 gnd OAI21X1_78/A OAI21X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1694 OAI21X1_79/a_2_6# OAI21X1_78/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1695 XNOR2X1_58/A OAI21X1_79/C OAI21X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1696 OAI21X1_78/a_9_54# OAI21X1_78/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1697 XOR2X1_82/A OAI21X1_78/B OAI21X1_78/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1698 vdd OAI21X1_78/C XOR2X1_82/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1699 gnd OAI21X1_78/A OAI21X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1700 OAI21X1_78/a_2_6# OAI21X1_78/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1701 XOR2X1_82/A OAI21X1_78/C OAI21X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1702 vdd XOR2X1_82/A XOR2X1_82/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1703 XOR2X1_82/a_18_54# XOR2X1_82/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1704 XOR2X1_82/Y XOR2X1_82/A XOR2X1_82/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1705 XOR2X1_82/a_35_54# XOR2X1_82/a_2_6# XOR2X1_82/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1706 vdd XOR2X1_82/B XOR2X1_82/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1707 XOR2X1_82/a_13_43# XOR2X1_82/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1708 gnd XOR2X1_82/A XOR2X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1709 XOR2X1_82/a_18_6# XOR2X1_82/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1710 XOR2X1_82/Y XOR2X1_82/a_2_6# XOR2X1_82/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1711 XOR2X1_82/a_35_6# XOR2X1_82/A XOR2X1_82/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1712 gnd XOR2X1_82/B XOR2X1_82/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1713 XOR2X1_82/a_13_43# XOR2X1_82/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1714 NOR2X1_43/a_9_54# AOI21X1_7/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1715 XOR2X1_85/B AOI21X1_7/B NOR2X1_43/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1716 XOR2X1_85/B AOI21X1_7/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1717 gnd AOI21X1_7/B XOR2X1_85/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 vdd AOI21X1_7/A AOI21X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M1719 AOI21X1_7/a_2_54# AOI21X1_7/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 INVX2_123/A XOR2X1_85/B AOI21X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1721 AOI21X1_7/a_12_6# AOI21X1_7/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1722 INVX2_123/A AOI21X1_7/B AOI21X1_7/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M1723 gnd XOR2X1_85/B INVX2_123/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1724 INVX2_123/Y INVX2_123/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1725 INVX2_123/Y INVX2_123/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1726 OAI22X1_18/a_9_54# INVX2_121/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1727 OAI22X1_18/Y INVX2_84/Y OAI22X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1728 OAI22X1_18/a_28_54# INVX2_99/Y OAI22X1_18/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1729 vdd XOR2X1_17/B OAI22X1_18/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1730 gnd INVX2_121/Y OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1731 OAI22X1_18/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1732 OAI22X1_18/Y INVX2_99/Y OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1733 OAI22X1_18/a_2_6# XOR2X1_17/B OAI22X1_18/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1734 OAI22X1_17/a_9_54# INVX2_122/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1735 OAI22X1_17/Y INVX2_84/Y OAI22X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1736 OAI22X1_17/a_28_54# INVX2_99/Y OAI22X1_17/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1737 vdd INVX2_87/Y OAI22X1_17/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1738 gnd INVX2_122/Y OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1739 OAI22X1_17/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1740 OAI22X1_17/Y INVX2_99/Y OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1741 OAI22X1_17/a_2_6# INVX2_87/Y OAI22X1_17/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1742 OAI22X1_16/a_9_54# INVX2_133/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1743 OAI22X1_16/Y INVX2_84/Y OAI22X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M1744 OAI22X1_16/a_28_54# INVX2_99/Y OAI22X1_16/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1745 vdd INVX2_17/Y OAI22X1_16/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1746 gnd INVX2_133/Y OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M1747 OAI22X1_16/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1748 OAI22X1_16/Y INVX2_99/Y OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1749 OAI22X1_16/a_2_6# INVX2_17/Y OAI22X1_16/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1750 INVX2_122/Y INVX2_122/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1751 INVX2_122/Y INVX2_122/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1752 INVX2_121/Y INVX2_121/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1753 INVX2_121/Y INVX2_121/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1754 vdd BUFX2_10/Y DFFPOSX1_87/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1755 DFFPOSX1_87/a_17_74# OAI21X1_76/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1756 DFFPOSX1_87/a_22_6# BUFX2_10/Y DFFPOSX1_87/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1757 DFFPOSX1_87/a_31_74# DFFPOSX1_87/a_2_6# DFFPOSX1_87/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1758 vdd DFFPOSX1_87/a_34_4# DFFPOSX1_87/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1759 DFFPOSX1_87/a_34_4# DFFPOSX1_87/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1760 DFFPOSX1_87/a_61_74# DFFPOSX1_87/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1761 DFFPOSX1_87/a_66_6# DFFPOSX1_87/a_2_6# DFFPOSX1_87/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1762 DFFPOSX1_87/a_76_84# BUFX2_10/Y DFFPOSX1_87/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1763 vdd out_MemBData[11] DFFPOSX1_87/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1764 gnd BUFX2_10/Y DFFPOSX1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1765 out_MemBData[11] DFFPOSX1_87/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1766 DFFPOSX1_87/a_17_6# OAI21X1_76/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1767 DFFPOSX1_87/a_22_6# DFFPOSX1_87/a_2_6# DFFPOSX1_87/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1768 DFFPOSX1_87/a_31_6# BUFX2_10/Y DFFPOSX1_87/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1769 gnd DFFPOSX1_87/a_34_4# DFFPOSX1_87/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1770 DFFPOSX1_87/a_34_4# DFFPOSX1_87/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1771 DFFPOSX1_87/a_61_6# DFFPOSX1_87/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1772 DFFPOSX1_87/a_66_6# BUFX2_10/Y DFFPOSX1_87/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1773 DFFPOSX1_87/a_76_6# DFFPOSX1_87/a_2_6# DFFPOSX1_87/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1774 gnd out_MemBData[11] DFFPOSX1_87/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1775 out_MemBData[11] DFFPOSX1_87/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1776 NOR2X1_41/a_9_54# INVX2_62/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1777 NOR2X1_41/Y NOR2X1_41/B NOR2X1_41/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1778 NOR2X1_41/Y INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1779 gnd NOR2X1_41/B NOR2X1_41/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1780 OAI21X1_77/a_9_54# NOR2X1_41/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1781 OAI21X1_76/C AND2X2_19/Y OAI21X1_77/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1782 vdd out_MemBData[11] OAI21X1_76/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1783 gnd NOR2X1_41/Y OAI21X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1784 OAI21X1_77/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1785 OAI21X1_76/C out_MemBData[11] OAI21X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1786 OAI21X1_76/a_9_54# INVX2_120/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1787 OAI21X1_76/Y OR2X2_0/Y OAI21X1_76/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1788 vdd OAI21X1_76/C OAI21X1_76/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1789 gnd INVX2_120/A OAI21X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1790 OAI21X1_76/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1791 OAI21X1_76/Y OAI21X1_76/C OAI21X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1792 NOR2X1_48/B INVX2_118/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1793 NOR2X1_48/B INVX2_118/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1794 vdd BUFX2_11/Y DFFPOSX1_85/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1795 DFFPOSX1_85/a_17_74# OAI21X1_83/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1796 DFFPOSX1_85/a_22_6# BUFX2_11/Y DFFPOSX1_85/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1797 DFFPOSX1_85/a_31_74# DFFPOSX1_85/a_2_6# DFFPOSX1_85/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1798 vdd DFFPOSX1_85/a_34_4# DFFPOSX1_85/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1799 DFFPOSX1_85/a_34_4# DFFPOSX1_85/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1800 DFFPOSX1_85/a_61_74# DFFPOSX1_85/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1801 DFFPOSX1_85/a_66_6# DFFPOSX1_85/a_2_6# DFFPOSX1_85/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1802 DFFPOSX1_85/a_76_84# BUFX2_11/Y DFFPOSX1_85/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1803 vdd out_MemBData[4] DFFPOSX1_85/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1804 gnd BUFX2_11/Y DFFPOSX1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1805 out_MemBData[4] DFFPOSX1_85/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1806 DFFPOSX1_85/a_17_6# OAI21X1_83/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1807 DFFPOSX1_85/a_22_6# DFFPOSX1_85/a_2_6# DFFPOSX1_85/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1808 DFFPOSX1_85/a_31_6# BUFX2_11/Y DFFPOSX1_85/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1809 gnd DFFPOSX1_85/a_34_4# DFFPOSX1_85/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1810 DFFPOSX1_85/a_34_4# DFFPOSX1_85/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1811 DFFPOSX1_85/a_61_6# DFFPOSX1_85/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1812 DFFPOSX1_85/a_66_6# BUFX2_11/Y DFFPOSX1_85/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1813 DFFPOSX1_85/a_76_6# DFFPOSX1_85/a_2_6# DFFPOSX1_85/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1814 gnd out_MemBData[4] DFFPOSX1_85/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1815 out_MemBData[4] DFFPOSX1_85/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1816 vdd BUFX2_11/Y DFFPOSX1_84/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1817 DFFPOSX1_84/a_17_74# OAI21X1_75/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1818 DFFPOSX1_84/a_22_6# BUFX2_11/Y DFFPOSX1_84/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1819 DFFPOSX1_84/a_31_74# DFFPOSX1_84/a_2_6# DFFPOSX1_84/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1820 vdd DFFPOSX1_84/a_34_4# DFFPOSX1_84/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1821 DFFPOSX1_84/a_34_4# DFFPOSX1_84/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1822 DFFPOSX1_84/a_61_74# DFFPOSX1_84/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1823 DFFPOSX1_84/a_66_6# DFFPOSX1_84/a_2_6# DFFPOSX1_84/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1824 DFFPOSX1_84/a_76_84# BUFX2_11/Y DFFPOSX1_84/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1825 vdd out_MemBData[5] DFFPOSX1_84/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1826 gnd BUFX2_11/Y DFFPOSX1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1827 out_MemBData[5] DFFPOSX1_84/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1828 DFFPOSX1_84/a_17_6# OAI21X1_75/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1829 DFFPOSX1_84/a_22_6# DFFPOSX1_84/a_2_6# DFFPOSX1_84/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1830 DFFPOSX1_84/a_31_6# BUFX2_11/Y DFFPOSX1_84/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1831 gnd DFFPOSX1_84/a_34_4# DFFPOSX1_84/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1832 DFFPOSX1_84/a_34_4# DFFPOSX1_84/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1833 DFFPOSX1_84/a_61_6# DFFPOSX1_84/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1834 DFFPOSX1_84/a_66_6# BUFX2_11/Y DFFPOSX1_84/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1835 DFFPOSX1_84/a_76_6# DFFPOSX1_84/a_2_6# DFFPOSX1_84/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1836 gnd out_MemBData[5] DFFPOSX1_84/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1837 out_MemBData[5] DFFPOSX1_84/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1838 OAI21X1_75/a_9_54# INVX2_117/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1839 OAI21X1_75/Y OR2X2_0/Y OAI21X1_75/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1840 vdd OAI21X1_81/Y OAI21X1_75/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1841 gnd INVX2_117/A OAI21X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1842 OAI21X1_75/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1843 OAI21X1_75/Y OAI21X1_81/Y OAI21X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1844 NOR2X1_46/B INVX2_117/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1845 NOR2X1_46/B INVX2_117/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1846 INVX2_116/Y INVX2_116/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1847 INVX2_116/Y INVX2_116/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1848 vdd con_count[2] AOI22X1_88/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1849 AOI22X1_88/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1850 INVX2_116/A INVX2_126/A AOI22X1_88/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1851 AOI22X1_88/a_2_54# AOI22X1_88/C INVX2_116/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1852 AOI22X1_88/a_11_6# con_count[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1853 INVX2_116/A INVX2_126/Y AOI22X1_88/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1854 AOI22X1_88/a_28_6# INVX2_126/A INVX2_116/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1855 gnd AOI22X1_88/C AOI22X1_88/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1856 vdd INVX2_43/Y DFFPOSX1_82/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1857 DFFPOSX1_82/a_17_74# INVX2_116/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1858 DFFPOSX1_82/a_22_6# INVX2_43/Y DFFPOSX1_82/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1859 DFFPOSX1_82/a_31_74# DFFPOSX1_82/a_2_6# DFFPOSX1_82/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1860 vdd DFFPOSX1_82/a_34_4# DFFPOSX1_82/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1861 DFFPOSX1_82/a_34_4# DFFPOSX1_82/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1862 DFFPOSX1_82/a_61_74# DFFPOSX1_82/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1863 DFFPOSX1_82/a_66_6# DFFPOSX1_82/a_2_6# DFFPOSX1_82/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1864 DFFPOSX1_82/a_76_84# INVX2_43/Y DFFPOSX1_82/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1865 vdd con_count[2] DFFPOSX1_82/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1866 gnd INVX2_43/Y DFFPOSX1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1867 con_count[2] DFFPOSX1_82/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1868 DFFPOSX1_82/a_17_6# INVX2_116/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1869 DFFPOSX1_82/a_22_6# DFFPOSX1_82/a_2_6# DFFPOSX1_82/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1870 DFFPOSX1_82/a_31_6# INVX2_43/Y DFFPOSX1_82/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1871 gnd DFFPOSX1_82/a_34_4# DFFPOSX1_82/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 DFFPOSX1_82/a_34_4# DFFPOSX1_82/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1873 DFFPOSX1_82/a_61_6# DFFPOSX1_82/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1874 DFFPOSX1_82/a_66_6# INVX2_43/Y DFFPOSX1_82/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1875 DFFPOSX1_82/a_76_6# DFFPOSX1_82/a_2_6# DFFPOSX1_82/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1876 gnd con_count[2] DFFPOSX1_82/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1877 con_count[2] DFFPOSX1_82/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1878 vdd con_count[3] HAX1_13/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1879 HAX1_13/a_2_74# HAX1_13/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1880 vdd HAX1_13/a_2_74# HAX1_12/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1881 HAX1_13/a_41_74# HAX1_13/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M1882 HAX1_13/a_49_54# HAX1_13/B HAX1_13/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1883 vdd con_count[3] HAX1_13/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1884 HAX1_13/YS HAX1_13/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1885 HAX1_13/a_9_6# con_count[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1886 HAX1_13/a_2_74# HAX1_13/B HAX1_13/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1887 gnd HAX1_13/a_2_74# HAX1_12/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1888 HAX1_13/a_38_6# HAX1_13/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M1889 HAX1_13/a_41_74# HAX1_13/B HAX1_13/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1890 HAX1_13/a_38_6# con_count[3] HAX1_13/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1891 HAX1_13/YS HAX1_13/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1892 NOR2X1_40/a_9_54# con_count[5] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1893 NOR2X1_40/Y con_count[4] NOR2X1_40/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1894 NOR2X1_40/Y con_count[5] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1895 gnd con_count[4] NOR2X1_40/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1896 vdd con_count[4] HAX1_12/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1897 HAX1_12/a_2_74# HAX1_12/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1898 vdd HAX1_12/a_2_74# HAX1_11/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1899 HAX1_12/a_41_74# HAX1_12/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M1900 HAX1_12/a_49_54# HAX1_12/B HAX1_12/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1901 vdd con_count[4] HAX1_12/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1902 HAX1_12/YS HAX1_12/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1903 HAX1_12/a_9_6# con_count[4] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1904 HAX1_12/a_2_74# HAX1_12/B HAX1_12/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1905 gnd HAX1_12/a_2_74# HAX1_11/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1906 HAX1_12/a_38_6# HAX1_12/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M1907 HAX1_12/a_41_74# HAX1_12/B HAX1_12/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1908 HAX1_12/a_38_6# con_count[4] HAX1_12/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1909 HAX1_12/YS HAX1_12/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1910 vdd con_count[5] AOI22X1_87/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1911 AOI22X1_87/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1912 INVX2_124/A INVX2_126/A AOI22X1_87/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1913 AOI22X1_87/a_2_54# AOI22X1_87/C INVX2_124/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1914 AOI22X1_87/a_11_6# con_count[5] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1915 INVX2_124/A INVX2_126/Y AOI22X1_87/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1916 AOI22X1_87/a_28_6# INVX2_126/A INVX2_124/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1917 gnd AOI22X1_87/C AOI22X1_87/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1918 vdd out_MuxData[4] XOR2X1_84/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1919 XOR2X1_84/a_18_54# XOR2X1_84/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1920 XOR2X1_83/B out_MuxData[4] XOR2X1_84/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1921 XOR2X1_84/a_35_54# XOR2X1_84/a_2_6# XOR2X1_83/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1922 vdd XOR2X1_84/B XOR2X1_84/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1923 XOR2X1_84/a_13_43# XOR2X1_84/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1924 gnd out_MuxData[4] XOR2X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1925 XOR2X1_84/a_18_6# XOR2X1_84/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1926 XOR2X1_83/B XOR2X1_84/a_2_6# XOR2X1_84/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1927 XOR2X1_84/a_35_6# out_MuxData[4] XOR2X1_83/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1928 gnd XOR2X1_84/B XOR2X1_84/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1929 XOR2X1_84/a_13_43# XOR2X1_84/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1930 vdd XOR2X1_83/B AOI22X1_92/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1931 AOI22X1_92/a_2_54# out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1932 NOR2X1_45/B out_MuxData[1] AOI22X1_92/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1933 AOI22X1_92/a_2_54# XOR2X1_83/Y NOR2X1_45/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1934 AOI22X1_92/a_11_6# XOR2X1_83/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1935 NOR2X1_45/B out_MuxData[2] AOI22X1_92/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1936 AOI22X1_92/a_28_6# out_MuxData[1] NOR2X1_45/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1937 gnd XOR2X1_83/Y AOI22X1_92/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1938 vdd out_MuxData[2] XOR2X1_83/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1939 XOR2X1_83/a_18_54# XOR2X1_83/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1940 XOR2X1_83/Y out_MuxData[2] XOR2X1_83/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1941 XOR2X1_83/a_35_54# XOR2X1_83/a_2_6# XOR2X1_83/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1942 vdd XOR2X1_83/B XOR2X1_83/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1943 XOR2X1_83/a_13_43# XOR2X1_83/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1944 gnd out_MuxData[2] XOR2X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1945 XOR2X1_83/a_18_6# XOR2X1_83/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1946 XOR2X1_83/Y XOR2X1_83/a_2_6# XOR2X1_83/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1947 XOR2X1_83/a_35_6# out_MuxData[2] XOR2X1_83/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1948 gnd XOR2X1_83/B XOR2X1_83/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1949 XOR2X1_83/a_13_43# XOR2X1_83/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1950 vdd XOR2X1_69/A XNOR2X1_55/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1951 XNOR2X1_55/a_18_54# XNOR2X1_55/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1952 XOR2X1_91/A XNOR2X1_55/a_2_6# XNOR2X1_55/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1953 XNOR2X1_55/a_35_54# XOR2X1_69/A XOR2X1_91/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1954 vdd XOR2X1_79/Y XNOR2X1_55/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1955 XNOR2X1_55/a_12_41# XOR2X1_79/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1956 gnd XOR2X1_69/A XNOR2X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1957 XNOR2X1_55/a_18_6# XNOR2X1_55/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1958 XOR2X1_91/A XOR2X1_69/A XNOR2X1_55/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1959 XNOR2X1_55/a_35_6# XNOR2X1_55/a_2_6# XOR2X1_91/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1960 gnd XOR2X1_79/Y XNOR2X1_55/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1961 XNOR2X1_55/a_12_41# XOR2X1_79/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1962 vdd OAI22X1_6/C XNOR2X1_54/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1963 XNOR2X1_54/a_18_54# XNOR2X1_54/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1964 AND2X2_40/A XNOR2X1_54/a_2_6# XNOR2X1_54/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1965 XNOR2X1_54/a_35_54# OAI22X1_6/C AND2X2_40/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1966 vdd XOR2X1_78/Y XNOR2X1_54/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1967 XNOR2X1_54/a_12_41# XOR2X1_78/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1968 gnd OAI22X1_6/C XNOR2X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1969 XNOR2X1_54/a_18_6# XNOR2X1_54/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1970 AND2X2_40/A OAI22X1_6/C XNOR2X1_54/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1971 XNOR2X1_54/a_35_6# XNOR2X1_54/a_2_6# AND2X2_40/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1972 gnd XOR2X1_78/Y XNOR2X1_54/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1973 XNOR2X1_54/a_12_41# XOR2X1_78/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1974 vdd NOR2X1_44/B XNOR2X1_53/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1975 XNOR2X1_53/a_18_54# XNOR2X1_53/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1976 OAI21X1_89/B XNOR2X1_53/a_2_6# XNOR2X1_53/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1977 XNOR2X1_53/a_35_54# NOR2X1_44/B OAI21X1_89/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1978 vdd NOR2X1_44/A XNOR2X1_53/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1979 XNOR2X1_53/a_12_41# NOR2X1_44/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1980 gnd NOR2X1_44/B XNOR2X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1981 XNOR2X1_53/a_18_6# XNOR2X1_53/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1982 OAI21X1_89/B NOR2X1_44/B XNOR2X1_53/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1983 XNOR2X1_53/a_35_6# XNOR2X1_53/a_2_6# OAI21X1_89/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1984 gnd NOR2X1_44/A XNOR2X1_53/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1985 XNOR2X1_53/a_12_41# NOR2X1_44/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1986 vdd XOR2X1_17/B XNOR2X1_52/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1987 XNOR2X1_52/a_18_54# XNOR2X1_52/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1988 XOR2X1_87/A XNOR2X1_52/a_2_6# XNOR2X1_52/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1989 XNOR2X1_52/a_35_54# XOR2X1_17/B XOR2X1_87/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1990 vdd XOR2X1_76/Y XNOR2X1_52/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1991 XNOR2X1_52/a_12_41# XOR2X1_76/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1992 gnd XOR2X1_17/B XNOR2X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1993 XNOR2X1_52/a_18_6# XNOR2X1_52/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1994 XOR2X1_87/A XOR2X1_17/B XNOR2X1_52/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1995 XNOR2X1_52/a_35_6# XNOR2X1_52/a_2_6# XOR2X1_87/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1996 gnd XOR2X1_76/Y XNOR2X1_52/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1997 XNOR2X1_52/a_12_41# XOR2X1_76/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1998 vdd out_MuxData[11] AOI22X1_90/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1999 AOI22X1_90/a_2_54# out_MuxData[8] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2000 NOR2X1_44/B out_MuxData[7] AOI22X1_90/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2001 AOI22X1_90/a_2_54# XOR2X1_77/Y NOR2X1_44/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2002 AOI22X1_90/a_11_6# out_MuxData[11] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2003 NOR2X1_44/B out_MuxData[8] AOI22X1_90/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2004 AOI22X1_90/a_28_6# out_MuxData[7] NOR2X1_44/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2005 gnd XOR2X1_77/Y AOI22X1_90/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2006 OAI21X1_79/C OAI21X1_78/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2007 vdd OAI21X1_78/B OAI21X1_79/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2008 NAND2X1_40/a_9_6# OAI21X1_78/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2009 OAI21X1_79/C OAI21X1_78/B NAND2X1_40/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2010 vdd NOR2X1_42/B XNOR2X1_51/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2011 XNOR2X1_51/a_18_54# XNOR2X1_51/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2012 OAI21X1_78/B XNOR2X1_51/a_2_6# XNOR2X1_51/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2013 XNOR2X1_51/a_35_54# NOR2X1_42/B OAI21X1_78/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2014 vdd NOR2X1_42/A XNOR2X1_51/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2015 XNOR2X1_51/a_12_41# NOR2X1_42/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2016 gnd NOR2X1_42/B XNOR2X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2017 XNOR2X1_51/a_18_6# XNOR2X1_51/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2018 OAI21X1_78/B NOR2X1_42/B XNOR2X1_51/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2019 XNOR2X1_51/a_35_6# XNOR2X1_51/a_2_6# OAI21X1_78/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2020 gnd NOR2X1_42/A XNOR2X1_51/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2021 XNOR2X1_51/a_12_41# NOR2X1_42/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2022 NOR2X1_42/a_9_54# NOR2X1_42/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2023 XOR2X1_82/B NOR2X1_42/B NOR2X1_42/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2024 XOR2X1_82/B NOR2X1_42/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2025 gnd NOR2X1_42/B XOR2X1_82/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2026 vdd XOR2X1_81/A XOR2X1_81/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2027 XOR2X1_81/a_18_54# XOR2X1_81/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2028 XOR2X1_81/Y XOR2X1_81/A XOR2X1_81/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2029 XOR2X1_81/a_35_54# XOR2X1_81/a_2_6# XOR2X1_81/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2030 vdd INVX2_17/Y XOR2X1_81/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2031 XOR2X1_81/a_13_43# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2032 gnd XOR2X1_81/A XOR2X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2033 XOR2X1_81/a_18_6# XOR2X1_81/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2034 XOR2X1_81/Y XOR2X1_81/a_2_6# XOR2X1_81/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2035 XOR2X1_81/a_35_6# XOR2X1_81/A XOR2X1_81/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2036 gnd INVX2_17/Y XOR2X1_81/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2037 XOR2X1_81/a_13_43# INVX2_17/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2038 vdd out_MuxData[7] AOI22X1_89/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2039 AOI22X1_89/a_2_54# out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2040 OAI21X1_87/A out_MuxData[11] AOI22X1_89/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2041 AOI22X1_89/a_2_54# XOR2X1_81/Y OAI21X1_87/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2042 AOI22X1_89/a_11_6# out_MuxData[7] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2043 OAI21X1_87/A out_MuxData[1] AOI22X1_89/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2044 AOI22X1_89/a_28_6# out_MuxData[11] OAI21X1_87/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2045 gnd XOR2X1_81/Y AOI22X1_89/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2046 vdd INVX2_87/Y XNOR2X1_50/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2047 XNOR2X1_50/a_18_54# XNOR2X1_50/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2048 AND2X2_36/B XNOR2X1_50/a_2_6# XNOR2X1_50/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2049 XNOR2X1_50/a_35_54# INVX2_87/Y AND2X2_36/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2050 vdd XOR2X1_81/Y XNOR2X1_50/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2051 XNOR2X1_50/a_12_41# XOR2X1_81/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2052 gnd INVX2_87/Y XNOR2X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2053 XNOR2X1_50/a_18_6# XNOR2X1_50/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2054 AND2X2_36/B INVX2_87/Y XNOR2X1_50/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2055 XNOR2X1_50/a_35_6# XNOR2X1_50/a_2_6# AND2X2_36/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2056 gnd XOR2X1_81/Y XNOR2X1_50/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2057 XNOR2X1_50/a_12_41# XOR2X1_81/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2058 vdd BUFX2_10/Y DFFPOSX1_89/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2059 DFFPOSX1_89/a_17_74# OAI22X1_18/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2060 DFFPOSX1_89/a_22_6# BUFX2_10/Y DFFPOSX1_89/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2061 DFFPOSX1_89/a_31_74# DFFPOSX1_89/a_2_6# DFFPOSX1_89/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2062 vdd DFFPOSX1_89/a_34_4# DFFPOSX1_89/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2063 DFFPOSX1_89/a_34_4# DFFPOSX1_89/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2064 DFFPOSX1_89/a_61_74# DFFPOSX1_89/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2065 DFFPOSX1_89/a_66_6# DFFPOSX1_89/a_2_6# DFFPOSX1_89/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2066 DFFPOSX1_89/a_76_84# BUFX2_10/Y DFFPOSX1_89/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2067 vdd out_MuxData[8] DFFPOSX1_89/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2068 gnd BUFX2_10/Y DFFPOSX1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2069 out_MuxData[8] DFFPOSX1_89/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2070 DFFPOSX1_89/a_17_6# OAI22X1_18/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2071 DFFPOSX1_89/a_22_6# DFFPOSX1_89/a_2_6# DFFPOSX1_89/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2072 DFFPOSX1_89/a_31_6# BUFX2_10/Y DFFPOSX1_89/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2073 gnd DFFPOSX1_89/a_34_4# DFFPOSX1_89/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2074 DFFPOSX1_89/a_34_4# DFFPOSX1_89/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2075 DFFPOSX1_89/a_61_6# DFFPOSX1_89/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2076 DFFPOSX1_89/a_66_6# BUFX2_10/Y DFFPOSX1_89/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2077 DFFPOSX1_89/a_76_6# DFFPOSX1_89/a_2_6# DFFPOSX1_89/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2078 gnd out_MuxData[8] DFFPOSX1_89/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2079 out_MuxData[8] DFFPOSX1_89/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2080 vdd INVX2_61/Y DFFPOSX1_88/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2081 DFFPOSX1_88/a_17_74# OAI22X1_15/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2082 DFFPOSX1_88/a_22_6# INVX2_61/Y DFFPOSX1_88/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2083 DFFPOSX1_88/a_31_74# DFFPOSX1_88/a_2_6# DFFPOSX1_88/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2084 vdd DFFPOSX1_88/a_34_4# DFFPOSX1_88/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2085 DFFPOSX1_88/a_34_4# DFFPOSX1_88/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2086 DFFPOSX1_88/a_61_74# DFFPOSX1_88/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2087 DFFPOSX1_88/a_66_6# DFFPOSX1_88/a_2_6# DFFPOSX1_88/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2088 DFFPOSX1_88/a_76_84# INVX2_61/Y DFFPOSX1_88/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2089 vdd INVX2_121/A DFFPOSX1_88/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2090 gnd INVX2_61/Y DFFPOSX1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2091 INVX2_121/A DFFPOSX1_88/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2092 DFFPOSX1_88/a_17_6# OAI22X1_15/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2093 DFFPOSX1_88/a_22_6# DFFPOSX1_88/a_2_6# DFFPOSX1_88/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2094 DFFPOSX1_88/a_31_6# INVX2_61/Y DFFPOSX1_88/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2095 gnd DFFPOSX1_88/a_34_4# DFFPOSX1_88/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2096 DFFPOSX1_88/a_34_4# DFFPOSX1_88/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2097 DFFPOSX1_88/a_61_6# DFFPOSX1_88/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2098 DFFPOSX1_88/a_66_6# INVX2_61/Y DFFPOSX1_88/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2099 DFFPOSX1_88/a_76_6# DFFPOSX1_88/a_2_6# DFFPOSX1_88/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2100 gnd INVX2_121/A DFFPOSX1_88/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2101 INVX2_121/A DFFPOSX1_88/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2102 OAI22X1_15/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2103 OAI22X1_15/Y INVX2_121/Y OAI22X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2104 OAI22X1_15/a_28_54# INVX2_119/Y OAI22X1_15/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2105 vdd INVX2_62/Y OAI22X1_15/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2106 gnd BUFX2_4/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2107 OAI22X1_15/a_2_6# INVX2_121/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2108 OAI22X1_15/Y INVX2_119/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2109 OAI22X1_15/a_2_6# INVX2_62/Y OAI22X1_15/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2110 NOR2X1_41/B INVX2_120/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2111 NOR2X1_41/B INVX2_120/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2112 vdd BUFX2_10/Y DFFPOSX1_86/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2113 DFFPOSX1_86/a_17_74# OAI21X1_73/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2114 DFFPOSX1_86/a_22_6# BUFX2_10/Y DFFPOSX1_86/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2115 DFFPOSX1_86/a_31_74# DFFPOSX1_86/a_2_6# DFFPOSX1_86/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2116 vdd DFFPOSX1_86/a_34_4# DFFPOSX1_86/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2117 DFFPOSX1_86/a_34_4# DFFPOSX1_86/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2118 DFFPOSX1_86/a_61_74# DFFPOSX1_86/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2119 DFFPOSX1_86/a_66_6# DFFPOSX1_86/a_2_6# DFFPOSX1_86/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2120 DFFPOSX1_86/a_76_84# BUFX2_10/Y DFFPOSX1_86/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2121 vdd out_MemBData[10] DFFPOSX1_86/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2122 gnd BUFX2_10/Y DFFPOSX1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2123 out_MemBData[10] DFFPOSX1_86/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2124 DFFPOSX1_86/a_17_6# OAI21X1_73/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2125 DFFPOSX1_86/a_22_6# DFFPOSX1_86/a_2_6# DFFPOSX1_86/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2126 DFFPOSX1_86/a_31_6# BUFX2_10/Y DFFPOSX1_86/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2127 gnd DFFPOSX1_86/a_34_4# DFFPOSX1_86/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2128 DFFPOSX1_86/a_34_4# DFFPOSX1_86/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2129 DFFPOSX1_86/a_61_6# DFFPOSX1_86/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2130 DFFPOSX1_86/a_66_6# BUFX2_10/Y DFFPOSX1_86/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2131 DFFPOSX1_86/a_76_6# DFFPOSX1_86/a_2_6# DFFPOSX1_86/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2132 gnd out_MemBData[10] DFFPOSX1_86/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2133 out_MemBData[10] DFFPOSX1_86/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2134 INVX2_119/Y out_MemBData[8] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2135 INVX2_119/Y out_MemBData[8] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2136 vdd BUFX2_10/Y DFFPOSX1_83/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2137 DFFPOSX1_83/a_17_74# OAI21X1_71/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2138 DFFPOSX1_83/a_22_6# BUFX2_10/Y DFFPOSX1_83/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2139 DFFPOSX1_83/a_31_74# DFFPOSX1_83/a_2_6# DFFPOSX1_83/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2140 vdd DFFPOSX1_83/a_34_4# DFFPOSX1_83/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2141 DFFPOSX1_83/a_34_4# DFFPOSX1_83/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2142 DFFPOSX1_83/a_61_74# DFFPOSX1_83/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2143 DFFPOSX1_83/a_66_6# DFFPOSX1_83/a_2_6# DFFPOSX1_83/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2144 DFFPOSX1_83/a_76_84# BUFX2_10/Y DFFPOSX1_83/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2145 vdd out_MemBData[8] DFFPOSX1_83/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2146 gnd BUFX2_10/Y DFFPOSX1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2147 out_MemBData[8] DFFPOSX1_83/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2148 DFFPOSX1_83/a_17_6# OAI21X1_71/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2149 DFFPOSX1_83/a_22_6# DFFPOSX1_83/a_2_6# DFFPOSX1_83/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2150 DFFPOSX1_83/a_31_6# BUFX2_10/Y DFFPOSX1_83/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2151 gnd DFFPOSX1_83/a_34_4# DFFPOSX1_83/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2152 DFFPOSX1_83/a_34_4# DFFPOSX1_83/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2153 DFFPOSX1_83/a_61_6# DFFPOSX1_83/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2154 DFFPOSX1_83/a_66_6# BUFX2_10/Y DFFPOSX1_83/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2155 DFFPOSX1_83/a_76_6# DFFPOSX1_83/a_2_6# DFFPOSX1_83/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2156 gnd out_MemBData[8] DFFPOSX1_83/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2157 out_MemBData[8] DFFPOSX1_83/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2158 INVX2_130/A NOR2X1_22/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2159 vdd NOR2X1_39/Y INVX2_130/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2160 NAND2X1_39/a_9_6# NOR2X1_22/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2161 INVX2_130/A NOR2X1_39/Y NAND2X1_39/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2162 INVX2_118/A NOR2X1_31/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2163 vdd NOR2X1_39/Y INVX2_118/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2164 NAND2X1_38/a_9_6# NOR2X1_31/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2165 INVX2_118/A NOR2X1_39/Y NAND2X1_38/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2166 INVX2_128/A NOR2X1_21/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2167 vdd NOR2X1_39/Y INVX2_128/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2168 NAND2X1_37/a_9_6# NOR2X1_21/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2169 INVX2_128/A NOR2X1_39/Y NAND2X1_37/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2170 INVX2_117/A NOR2X1_30/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2171 vdd NOR2X1_39/Y INVX2_117/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2172 NAND2X1_36/a_9_6# NOR2X1_30/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2173 INVX2_117/A NOR2X1_39/Y NAND2X1_36/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2174 NOR2X1_39/a_9_54# NOR2X1_39/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2175 NOR2X1_39/Y con_count[3] NOR2X1_39/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2176 NOR2X1_39/Y NOR2X1_39/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2177 gnd con_count[3] NOR2X1_39/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2178 NOR2X1_39/A con_count[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2179 NOR2X1_39/A con_count[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2180 vdd BUFX2_9/Y DFFPOSX1_81/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2181 DFFPOSX1_81/a_17_74# AND2X2_33/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2182 DFFPOSX1_81/a_22_6# BUFX2_9/Y DFFPOSX1_81/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2183 DFFPOSX1_81/a_31_74# DFFPOSX1_81/a_2_6# DFFPOSX1_81/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2184 vdd DFFPOSX1_81/a_34_4# DFFPOSX1_81/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2185 DFFPOSX1_81/a_34_4# DFFPOSX1_81/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2186 DFFPOSX1_81/a_61_74# DFFPOSX1_81/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2187 DFFPOSX1_81/a_66_6# DFFPOSX1_81/a_2_6# DFFPOSX1_81/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2188 DFFPOSX1_81/a_76_84# BUFX2_9/Y DFFPOSX1_81/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2189 vdd AOI22X1_88/C DFFPOSX1_81/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2190 gnd BUFX2_9/Y DFFPOSX1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2191 AOI22X1_88/C DFFPOSX1_81/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2192 DFFPOSX1_81/a_17_6# AND2X2_33/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2193 DFFPOSX1_81/a_22_6# DFFPOSX1_81/a_2_6# DFFPOSX1_81/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2194 DFFPOSX1_81/a_31_6# BUFX2_9/Y DFFPOSX1_81/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2195 gnd DFFPOSX1_81/a_34_4# DFFPOSX1_81/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2196 DFFPOSX1_81/a_34_4# DFFPOSX1_81/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2197 DFFPOSX1_81/a_61_6# DFFPOSX1_81/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2198 DFFPOSX1_81/a_66_6# BUFX2_9/Y DFFPOSX1_81/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2199 DFFPOSX1_81/a_76_6# DFFPOSX1_81/a_2_6# DFFPOSX1_81/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2200 gnd AOI22X1_88/C DFFPOSX1_81/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2201 AOI22X1_88/C DFFPOSX1_81/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2202 AND2X2_33/a_2_6# HAX1_10/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2203 vdd INVX2_72/Y AND2X2_33/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2204 AND2X2_33/Y AND2X2_33/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2205 AND2X2_33/a_9_6# HAX1_10/YS AND2X2_33/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M2206 gnd INVX2_72/Y AND2X2_33/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2207 AND2X2_33/Y AND2X2_33/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2208 AND2X2_32/a_2_6# HAX1_11/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2209 vdd INVX2_72/Y AND2X2_32/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2210 AND2X2_32/Y AND2X2_32/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2211 AND2X2_32/a_9_6# HAX1_11/YS AND2X2_32/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M2212 gnd INVX2_72/Y AND2X2_32/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2213 AND2X2_32/Y AND2X2_32/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2214 vdd con_count[5] HAX1_11/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M2215 HAX1_11/a_2_74# HAX1_11/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2216 vdd HAX1_11/a_2_74# HAX1_9/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2217 HAX1_11/a_41_74# HAX1_11/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M2218 HAX1_11/a_49_54# HAX1_11/B HAX1_11/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2219 vdd con_count[5] HAX1_11/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2220 HAX1_11/YS HAX1_11/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2221 HAX1_11/a_9_6# con_count[5] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2222 HAX1_11/a_2_74# HAX1_11/B HAX1_11/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2223 gnd HAX1_11/a_2_74# HAX1_9/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M2224 HAX1_11/a_38_6# HAX1_11/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M2225 HAX1_11/a_41_74# HAX1_11/B HAX1_11/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2226 HAX1_11/a_38_6# con_count[5] HAX1_11/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2227 HAX1_11/YS HAX1_11/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2228 vdd BUFX2_9/Y DFFPOSX1_80/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2229 DFFPOSX1_80/a_17_74# AND2X2_32/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2230 DFFPOSX1_80/a_22_6# BUFX2_9/Y DFFPOSX1_80/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2231 DFFPOSX1_80/a_31_74# DFFPOSX1_80/a_2_6# DFFPOSX1_80/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2232 vdd DFFPOSX1_80/a_34_4# DFFPOSX1_80/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2233 DFFPOSX1_80/a_34_4# DFFPOSX1_80/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2234 DFFPOSX1_80/a_61_74# DFFPOSX1_80/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2235 DFFPOSX1_80/a_66_6# DFFPOSX1_80/a_2_6# DFFPOSX1_80/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2236 DFFPOSX1_80/a_76_84# BUFX2_9/Y DFFPOSX1_80/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2237 vdd AOI22X1_87/C DFFPOSX1_80/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2238 gnd BUFX2_9/Y DFFPOSX1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2239 AOI22X1_87/C DFFPOSX1_80/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2240 DFFPOSX1_80/a_17_6# AND2X2_32/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2241 DFFPOSX1_80/a_22_6# DFFPOSX1_80/a_2_6# DFFPOSX1_80/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2242 DFFPOSX1_80/a_31_6# BUFX2_9/Y DFFPOSX1_80/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2243 gnd DFFPOSX1_80/a_34_4# DFFPOSX1_80/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2244 DFFPOSX1_80/a_34_4# DFFPOSX1_80/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2245 DFFPOSX1_80/a_61_6# DFFPOSX1_80/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2246 DFFPOSX1_80/a_66_6# BUFX2_9/Y DFFPOSX1_80/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2247 DFFPOSX1_80/a_76_6# DFFPOSX1_80/a_2_6# DFFPOSX1_80/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2248 gnd AOI22X1_87/C DFFPOSX1_80/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2249 AOI22X1_87/C DFFPOSX1_80/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2250 XOR2X1_81/A out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2251 XOR2X1_81/A out_MuxData[1] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2252 vdd OAI22X1_6/C XOR2X1_79/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2253 XOR2X1_79/a_18_54# XOR2X1_79/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2254 XOR2X1_79/Y OAI22X1_6/C XOR2X1_79/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2255 XOR2X1_79/a_35_54# XOR2X1_79/a_2_6# XOR2X1_79/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2256 vdd INVX2_16/Y XOR2X1_79/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2257 XOR2X1_79/a_13_43# INVX2_16/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2258 gnd OAI22X1_6/C XOR2X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2259 XOR2X1_79/a_18_6# XOR2X1_79/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2260 XOR2X1_79/Y XOR2X1_79/a_2_6# XOR2X1_79/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2261 XOR2X1_79/a_35_6# OAI22X1_6/C XOR2X1_79/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2262 gnd INVX2_16/Y XOR2X1_79/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2263 XOR2X1_79/a_13_43# INVX2_16/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2264 vdd out_MuxData[6] AOI22X1_85/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2265 AOI22X1_85/a_2_54# out_MuxData[0] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2266 OAI21X1_91/A out_MuxData[10] AOI22X1_85/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2267 AOI22X1_85/a_2_54# XOR2X1_79/Y OAI21X1_91/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2268 AOI22X1_85/a_11_6# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2269 OAI21X1_91/A out_MuxData[0] AOI22X1_85/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2270 AOI22X1_85/a_28_6# out_MuxData[10] OAI21X1_91/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2271 gnd XOR2X1_79/Y AOI22X1_85/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2272 vdd out_MuxData[1] XOR2X1_78/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2273 XOR2X1_78/a_18_54# XOR2X1_78/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2274 XOR2X1_78/Y out_MuxData[1] XOR2X1_78/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2275 XOR2X1_78/a_35_54# XOR2X1_78/a_2_6# XOR2X1_78/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2276 vdd XOR2X1_78/B XOR2X1_78/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2277 XOR2X1_78/a_13_43# XOR2X1_78/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2278 gnd out_MuxData[1] XOR2X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2279 XOR2X1_78/a_18_6# XOR2X1_78/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2280 XOR2X1_78/Y XOR2X1_78/a_2_6# XOR2X1_78/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2281 XOR2X1_78/a_35_6# out_MuxData[1] XOR2X1_78/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2282 gnd XOR2X1_78/B XOR2X1_78/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2283 XOR2X1_78/a_13_43# XOR2X1_78/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2284 vdd XOR2X1_78/B AOI22X1_84/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2285 AOI22X1_84/a_2_54# out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2286 NOR2X1_44/A out_MuxData[0] AOI22X1_84/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2287 AOI22X1_84/a_2_54# XOR2X1_78/Y NOR2X1_44/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2288 AOI22X1_84/a_11_6# XOR2X1_78/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2289 NOR2X1_44/A out_MuxData[1] AOI22X1_84/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2290 AOI22X1_84/a_28_6# out_MuxData[0] NOR2X1_44/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2291 gnd XOR2X1_78/Y AOI22X1_84/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2292 vdd INVX2_87/Y XOR2X1_77/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2293 XOR2X1_77/a_18_54# XOR2X1_77/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2294 XOR2X1_77/Y INVX2_87/Y XOR2X1_77/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2295 XOR2X1_77/a_35_54# XOR2X1_77/a_2_6# XOR2X1_77/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2296 vdd XOR2X1_17/B XOR2X1_77/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2297 XOR2X1_77/a_13_43# XOR2X1_17/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2298 gnd INVX2_87/Y XOR2X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2299 XOR2X1_77/a_18_6# XOR2X1_77/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2300 XOR2X1_77/Y XOR2X1_77/a_2_6# XOR2X1_77/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2301 XOR2X1_77/a_35_6# INVX2_87/Y XOR2X1_77/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2302 gnd XOR2X1_17/B XOR2X1_77/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2303 XOR2X1_77/a_13_43# XOR2X1_17/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2304 vdd INVX2_17/Y XNOR2X1_48/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2305 XNOR2X1_48/a_18_54# XNOR2X1_48/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2306 XOR2X1_78/B XNOR2X1_48/a_2_6# XNOR2X1_48/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2307 XNOR2X1_48/a_35_54# INVX2_17/Y XOR2X1_78/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2308 vdd XOR2X1_77/Y XNOR2X1_48/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2309 XNOR2X1_48/a_12_41# XOR2X1_77/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2310 gnd INVX2_17/Y XNOR2X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2311 XNOR2X1_48/a_18_6# XNOR2X1_48/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2312 XOR2X1_78/B INVX2_17/Y XNOR2X1_48/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2313 XNOR2X1_48/a_35_6# XNOR2X1_48/a_2_6# XOR2X1_78/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2314 gnd XOR2X1_77/Y XNOR2X1_48/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2315 XNOR2X1_48/a_12_41# XOR2X1_77/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2316 vdd out_MuxData[4] AOI22X1_83/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2317 AOI22X1_83/a_2_54# out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2318 OAI21X1_78/A out_MuxData[8] AOI22X1_83/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2319 AOI22X1_83/a_2_54# XOR2X1_76/Y OAI21X1_78/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2320 AOI22X1_83/a_11_6# out_MuxData[4] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2321 OAI21X1_78/A out_MuxData[2] AOI22X1_83/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2322 AOI22X1_83/a_28_6# out_MuxData[8] OAI21X1_78/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2323 gnd XOR2X1_76/Y AOI22X1_83/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2324 vdd XOR2X1_75/Y AOI22X1_82/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2325 AOI22X1_82/a_2_54# out_MuxData[6] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2326 NOR2X1_42/B out_MuxData[11] AOI22X1_82/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2327 AOI22X1_82/a_2_54# out_MuxData[10] NOR2X1_42/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2328 AOI22X1_82/a_11_6# XOR2X1_75/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2329 NOR2X1_42/B out_MuxData[6] AOI22X1_82/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2330 AOI22X1_82/a_28_6# out_MuxData[11] NOR2X1_42/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2331 gnd out_MuxData[10] AOI22X1_82/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2332 OAI22X1_14/a_9_54# INVX2_134/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2333 OAI22X1_14/Y INVX2_84/Y OAI22X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2334 OAI22X1_14/a_28_54# INVX2_99/Y OAI22X1_14/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2335 vdd INVX2_16/Y OAI22X1_14/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2336 gnd INVX2_134/Y OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2337 OAI22X1_14/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2338 OAI22X1_14/Y INVX2_99/Y OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2339 OAI22X1_14/a_2_6# INVX2_16/Y OAI22X1_14/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2340 vdd BUFX2_11/Y DFFPOSX1_78/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2341 DFFPOSX1_78/a_17_74# OAI22X1_16/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2342 DFFPOSX1_78/a_22_6# BUFX2_11/Y DFFPOSX1_78/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2343 DFFPOSX1_78/a_31_74# DFFPOSX1_78/a_2_6# DFFPOSX1_78/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2344 vdd DFFPOSX1_78/a_34_4# DFFPOSX1_78/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2345 DFFPOSX1_78/a_34_4# DFFPOSX1_78/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2346 DFFPOSX1_78/a_61_74# DFFPOSX1_78/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2347 DFFPOSX1_78/a_66_6# DFFPOSX1_78/a_2_6# DFFPOSX1_78/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2348 DFFPOSX1_78/a_76_84# BUFX2_11/Y DFFPOSX1_78/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2349 vdd out_MuxData[7] DFFPOSX1_78/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2350 gnd BUFX2_11/Y DFFPOSX1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2351 out_MuxData[7] DFFPOSX1_78/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2352 DFFPOSX1_78/a_17_6# OAI22X1_16/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2353 DFFPOSX1_78/a_22_6# DFFPOSX1_78/a_2_6# DFFPOSX1_78/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2354 DFFPOSX1_78/a_31_6# BUFX2_11/Y DFFPOSX1_78/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2355 gnd DFFPOSX1_78/a_34_4# DFFPOSX1_78/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2356 DFFPOSX1_78/a_34_4# DFFPOSX1_78/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2357 DFFPOSX1_78/a_61_6# DFFPOSX1_78/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2358 DFFPOSX1_78/a_66_6# BUFX2_11/Y DFFPOSX1_78/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2359 DFFPOSX1_78/a_76_6# DFFPOSX1_78/a_2_6# DFFPOSX1_78/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2360 gnd out_MuxData[7] DFFPOSX1_78/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2361 out_MuxData[7] DFFPOSX1_78/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2362 INVX2_110/Y INVX2_110/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2363 INVX2_110/Y INVX2_110/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2364 vdd INVX2_61/Y DFFPOSX1_77/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2365 DFFPOSX1_77/a_17_74# OAI22X1_11/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2366 DFFPOSX1_77/a_22_6# INVX2_61/Y DFFPOSX1_77/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2367 DFFPOSX1_77/a_31_74# DFFPOSX1_77/a_2_6# DFFPOSX1_77/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2368 vdd DFFPOSX1_77/a_34_4# DFFPOSX1_77/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2369 DFFPOSX1_77/a_34_4# DFFPOSX1_77/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2370 DFFPOSX1_77/a_61_74# DFFPOSX1_77/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2371 DFFPOSX1_77/a_66_6# DFFPOSX1_77/a_2_6# DFFPOSX1_77/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2372 DFFPOSX1_77/a_76_84# INVX2_61/Y DFFPOSX1_77/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2373 vdd INVX2_110/A DFFPOSX1_77/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2374 gnd INVX2_61/Y DFFPOSX1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2375 INVX2_110/A DFFPOSX1_77/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2376 DFFPOSX1_77/a_17_6# OAI22X1_11/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2377 DFFPOSX1_77/a_22_6# DFFPOSX1_77/a_2_6# DFFPOSX1_77/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2378 DFFPOSX1_77/a_31_6# INVX2_61/Y DFFPOSX1_77/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2379 gnd DFFPOSX1_77/a_34_4# DFFPOSX1_77/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2380 DFFPOSX1_77/a_34_4# DFFPOSX1_77/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2381 DFFPOSX1_77/a_61_6# DFFPOSX1_77/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2382 DFFPOSX1_77/a_66_6# INVX2_61/Y DFFPOSX1_77/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2383 DFFPOSX1_77/a_76_6# DFFPOSX1_77/a_2_6# DFFPOSX1_77/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2384 gnd INVX2_110/A DFFPOSX1_77/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2385 INVX2_110/A DFFPOSX1_77/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2386 OAI22X1_11/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2387 OAI22X1_11/Y INVX2_110/Y OAI22X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2388 OAI22X1_11/a_28_54# INVX2_108/Y OAI22X1_11/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2389 vdd INVX2_62/Y OAI22X1_11/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2390 gnd BUFX2_4/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2391 OAI22X1_11/a_2_6# INVX2_110/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2392 OAI22X1_11/Y INVX2_108/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2393 OAI22X1_11/a_2_6# INVX2_62/Y OAI22X1_11/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2394 INVX2_108/Y out_MemBData[10] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2395 INVX2_108/Y out_MemBData[10] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2396 OAI21X1_74/a_9_54# NOR2X1_38/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2397 OAI21X1_73/C AND2X2_19/Y OAI21X1_74/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2398 vdd out_MemBData[10] OAI21X1_73/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2399 gnd NOR2X1_38/Y OAI21X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2400 OAI21X1_74/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2401 OAI21X1_73/C out_MemBData[10] OAI21X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2402 OAI21X1_73/a_9_54# INVX2_106/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2403 OAI21X1_73/Y OR2X2_0/Y OAI21X1_73/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2404 vdd OAI21X1_73/C OAI21X1_73/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2405 gnd INVX2_106/A OAI21X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2406 OAI21X1_73/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2407 OAI21X1_73/Y OAI21X1_73/C OAI21X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2408 NOR2X1_37/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2409 NOR2X1_37/Y INVX2_104/Y NOR2X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2410 NOR2X1_37/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2411 gnd INVX2_104/Y NOR2X1_37/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2412 OAI21X1_72/a_9_54# NOR2X1_37/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2413 OAI21X1_71/C AND2X2_19/Y OAI21X1_72/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2414 vdd out_MemBData[8] OAI21X1_71/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2415 gnd NOR2X1_37/Y OAI21X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2416 OAI21X1_72/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2417 OAI21X1_71/C out_MemBData[8] OAI21X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2418 OAI21X1_71/a_9_54# INVX2_104/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2419 OAI21X1_71/Y OR2X2_0/Y OAI21X1_71/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2420 vdd OAI21X1_71/C OAI21X1_71/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2421 gnd INVX2_104/A OAI21X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2422 OAI21X1_71/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2423 OAI21X1_71/Y OAI21X1_71/C OAI21X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2424 INVX2_104/Y INVX2_104/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2425 INVX2_104/Y INVX2_104/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2426 INVX2_120/A NOR2X1_36/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2427 vdd NOR2X1_22/Y INVX2_120/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2428 NAND2X1_35/a_9_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2429 INVX2_120/A NOR2X1_22/Y NAND2X1_35/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2430 INVX2_104/A NOR2X1_36/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2431 vdd NOR2X1_31/Y INVX2_104/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2432 NAND2X1_34/a_9_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2433 INVX2_104/A NOR2X1_31/Y NAND2X1_34/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2434 NOR2X1_36/a_9_54# INVX2_103/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2435 NOR2X1_36/Y con_count[2] NOR2X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2436 NOR2X1_36/Y INVX2_103/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2437 gnd con_count[2] NOR2X1_36/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2438 NOR2X1_35/a_9_54# INVX2_103/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2439 NOR2X1_35/Y NOR2X1_39/A NOR2X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2440 NOR2X1_35/Y INVX2_103/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2441 gnd NOR2X1_39/A NOR2X1_35/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2442 INVX2_103/Y con_count[3] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2443 INVX2_103/Y con_count[3] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2444 NAND3X1_29/Y con_count[3] vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M2445 vdd con_count[2] NAND3X1_29/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2446 NAND3X1_29/Y AND2X2_30/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2447 NAND3X1_29/a_9_6# con_count[3] gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2448 NAND3X1_29/a_14_6# con_count[2] NAND3X1_29/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2449 NAND3X1_29/Y AND2X2_30/Y NAND3X1_29/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M2450 vdd con_count[2] HAX1_10/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M2451 HAX1_10/a_2_74# HAX1_10/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2452 vdd HAX1_10/a_2_74# HAX1_13/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2453 HAX1_10/a_41_74# HAX1_10/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M2454 HAX1_10/a_49_54# HAX1_10/B HAX1_10/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2455 vdd con_count[2] HAX1_10/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2456 HAX1_10/YS HAX1_10/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2457 HAX1_10/a_9_6# con_count[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2458 HAX1_10/a_2_74# HAX1_10/B HAX1_10/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2459 gnd HAX1_10/a_2_74# HAX1_13/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M2460 HAX1_10/a_38_6# HAX1_10/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M2461 HAX1_10/a_41_74# HAX1_10/B HAX1_10/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2462 HAX1_10/a_38_6# con_count[2] HAX1_10/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2463 HAX1_10/YS HAX1_10/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2464 AND2X2_31/a_2_6# HAX1_9/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2465 vdd INVX2_72/Y AND2X2_31/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2466 AND2X2_31/Y AND2X2_31/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2467 AND2X2_31/a_9_6# HAX1_9/YS AND2X2_31/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M2468 gnd INVX2_72/Y AND2X2_31/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2469 AND2X2_31/Y AND2X2_31/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2470 vdd con_count[6] HAX1_9/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M2471 HAX1_9/a_2_74# HAX1_9/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2472 vdd HAX1_9/a_2_74# HAX1_7/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2473 HAX1_9/a_41_74# HAX1_9/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M2474 HAX1_9/a_49_54# HAX1_9/B HAX1_9/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2475 vdd con_count[6] HAX1_9/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2476 HAX1_9/YS HAX1_9/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2477 HAX1_9/a_9_6# con_count[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2478 HAX1_9/a_2_74# HAX1_9/B HAX1_9/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2479 gnd HAX1_9/a_2_74# HAX1_7/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M2480 HAX1_9/a_38_6# HAX1_9/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M2481 HAX1_9/a_41_74# HAX1_9/B HAX1_9/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2482 HAX1_9/a_38_6# con_count[6] HAX1_9/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2483 HAX1_9/YS HAX1_9/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2484 vdd BUFX2_9/Y DFFPOSX1_73/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2485 DFFPOSX1_73/a_17_74# AND2X2_31/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2486 DFFPOSX1_73/a_22_6# BUFX2_9/Y DFFPOSX1_73/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2487 DFFPOSX1_73/a_31_74# DFFPOSX1_73/a_2_6# DFFPOSX1_73/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2488 vdd DFFPOSX1_73/a_34_4# DFFPOSX1_73/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2489 DFFPOSX1_73/a_34_4# DFFPOSX1_73/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2490 DFFPOSX1_73/a_61_74# DFFPOSX1_73/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2491 DFFPOSX1_73/a_66_6# DFFPOSX1_73/a_2_6# DFFPOSX1_73/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2492 DFFPOSX1_73/a_76_84# BUFX2_9/Y DFFPOSX1_73/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2493 vdd AOI22X1_79/C DFFPOSX1_73/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2494 gnd BUFX2_9/Y DFFPOSX1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2495 AOI22X1_79/C DFFPOSX1_73/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2496 DFFPOSX1_73/a_17_6# AND2X2_31/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2497 DFFPOSX1_73/a_22_6# DFFPOSX1_73/a_2_6# DFFPOSX1_73/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2498 DFFPOSX1_73/a_31_6# BUFX2_9/Y DFFPOSX1_73/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2499 gnd DFFPOSX1_73/a_34_4# DFFPOSX1_73/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2500 DFFPOSX1_73/a_34_4# DFFPOSX1_73/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2501 DFFPOSX1_73/a_61_6# DFFPOSX1_73/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2502 DFFPOSX1_73/a_66_6# BUFX2_9/Y DFFPOSX1_73/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2503 DFFPOSX1_73/a_76_6# DFFPOSX1_73/a_2_6# DFFPOSX1_73/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2504 gnd AOI22X1_79/C DFFPOSX1_73/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2505 AOI22X1_79/C DFFPOSX1_73/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2506 vdd con_count[6] AOI22X1_79/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2507 AOI22X1_79/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2508 INVX2_102/A INVX2_126/A AOI22X1_79/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2509 AOI22X1_79/a_2_54# AOI22X1_79/C INVX2_102/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2510 AOI22X1_79/a_11_6# con_count[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2511 INVX2_102/A INVX2_126/Y AOI22X1_79/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2512 AOI22X1_79/a_28_6# INVX2_126/A INVX2_102/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2513 gnd AOI22X1_79/C AOI22X1_79/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2514 vdd out_MuxData[8] AOI22X1_86/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2515 AOI22X1_86/a_2_54# out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2516 NOR2X1_45/A out_MuxData[4] AOI22X1_86/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2517 AOI22X1_86/a_2_54# XOR2X1_84/B NOR2X1_45/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2518 AOI22X1_86/a_11_6# out_MuxData[8] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2519 NOR2X1_45/A out_MuxData[9] AOI22X1_86/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2520 AOI22X1_86/a_28_6# out_MuxData[4] NOR2X1_45/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2521 gnd XOR2X1_84/B AOI22X1_86/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2522 vdd XOR2X1_17/B XOR2X1_80/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2523 XOR2X1_80/a_18_54# XOR2X1_80/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2524 XOR2X1_84/B XOR2X1_17/B XOR2X1_80/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2525 XOR2X1_80/a_35_54# XOR2X1_80/a_2_6# XOR2X1_84/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2526 vdd XOR2X1_69/B XOR2X1_80/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2527 XOR2X1_80/a_13_43# XOR2X1_69/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2528 gnd XOR2X1_17/B XOR2X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2529 XOR2X1_80/a_18_6# XOR2X1_80/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2530 XOR2X1_84/B XOR2X1_80/a_2_6# XOR2X1_80/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2531 XOR2X1_80/a_35_6# XOR2X1_17/B XOR2X1_84/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2532 gnd XOR2X1_69/B XOR2X1_80/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2533 XOR2X1_80/a_13_43# XOR2X1_69/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2534 XOR2X1_69/B out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2535 XOR2X1_69/B out_MuxData[9] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2536 XOR2X1_17/B out_MuxData[8] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2537 XOR2X1_17/B out_MuxData[8] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2538 XOR2X1_69/A out_MuxData[10] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2539 XOR2X1_69/A out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2540 vdd XOR2X1_69/B XNOR2X1_49/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2541 XNOR2X1_49/a_18_54# XNOR2X1_49/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2542 XOR2X1_90/A XNOR2X1_49/a_2_6# XNOR2X1_49/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2543 XNOR2X1_49/a_35_54# XOR2X1_69/B XOR2X1_90/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2544 vdd XOR2X1_71/Y XNOR2X1_49/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2545 XNOR2X1_49/a_12_41# XOR2X1_71/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2546 gnd XOR2X1_69/B XNOR2X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2547 XNOR2X1_49/a_18_6# XNOR2X1_49/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2548 XOR2X1_90/A XOR2X1_69/B XNOR2X1_49/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2549 XNOR2X1_49/a_35_6# XNOR2X1_49/a_2_6# XOR2X1_90/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2550 gnd XOR2X1_71/Y XNOR2X1_49/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2551 XNOR2X1_49/a_12_41# XOR2X1_71/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2552 NOR2X1_16/B AOI22X1_99/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M2553 vdd AOI22X1_96/Y NOR2X1_16/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2554 NOR2X1_16/B AND2X2_17/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2555 NAND3X1_30/a_9_6# AOI22X1_99/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2556 NAND3X1_30/a_14_6# AOI22X1_96/Y NAND3X1_30/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2557 NOR2X1_16/B AND2X2_17/Y NAND3X1_30/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M2558 vdd out_MuxData[4] XOR2X1_76/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2559 XOR2X1_76/a_18_54# XOR2X1_76/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2560 XOR2X1_76/Y out_MuxData[4] XOR2X1_76/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2561 XOR2X1_76/a_35_54# XOR2X1_76/a_2_6# XOR2X1_76/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2562 vdd out_MuxData[2] XOR2X1_76/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2563 XOR2X1_76/a_13_43# out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2564 gnd out_MuxData[4] XOR2X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2565 XOR2X1_76/a_18_6# XOR2X1_76/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2566 XOR2X1_76/Y XOR2X1_76/a_2_6# XOR2X1_76/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2567 XOR2X1_76/a_35_6# out_MuxData[4] XOR2X1_76/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2568 gnd out_MuxData[2] XOR2X1_76/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2569 XOR2X1_76/a_13_43# out_MuxData[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2570 vdd XOR2X1_69/A XOR2X1_75/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2571 XOR2X1_75/a_18_54# XOR2X1_75/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2572 XOR2X1_75/Y XOR2X1_69/A XOR2X1_75/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2573 XOR2X1_75/a_35_54# XOR2X1_75/a_2_6# XOR2X1_75/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2574 vdd INVX2_87/Y XOR2X1_75/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2575 XOR2X1_75/a_13_43# INVX2_87/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2576 gnd XOR2X1_69/A XOR2X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2577 XOR2X1_75/a_18_6# XOR2X1_75/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2578 XOR2X1_75/Y XOR2X1_75/a_2_6# XOR2X1_75/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2579 XOR2X1_75/a_35_6# XOR2X1_69/A XOR2X1_75/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2580 gnd INVX2_87/Y XOR2X1_75/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2581 XOR2X1_75/a_13_43# INVX2_87/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2582 vdd INVX2_16/Y XNOR2X1_47/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2583 XNOR2X1_47/a_18_54# XNOR2X1_47/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2584 XOR2X1_70/B XNOR2X1_47/a_2_6# XNOR2X1_47/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2585 XNOR2X1_47/a_35_54# INVX2_16/Y XOR2X1_70/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2586 vdd XOR2X1_75/Y XNOR2X1_47/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2587 XNOR2X1_47/a_12_41# XOR2X1_75/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2588 gnd INVX2_16/Y XNOR2X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2589 XNOR2X1_47/a_18_6# XNOR2X1_47/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2590 XOR2X1_70/B INVX2_16/Y XNOR2X1_47/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2591 XNOR2X1_47/a_35_6# XNOR2X1_47/a_2_6# XOR2X1_70/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2592 gnd XOR2X1_75/Y XNOR2X1_47/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2593 XNOR2X1_47/a_12_41# XOR2X1_75/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2594 vdd out_MuxData[10] AOI22X1_81/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2595 AOI22X1_81/a_2_54# out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2596 AOI21X1_7/A out_MuxData[5] AOI22X1_81/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2597 AOI22X1_81/a_2_54# XOR2X1_68/B AOI21X1_7/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2598 AOI22X1_81/a_11_6# out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2599 AOI21X1_7/A out_MuxData[9] AOI22X1_81/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2600 AOI22X1_81/a_28_6# out_MuxData[5] AOI21X1_7/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2601 gnd XOR2X1_68/B AOI22X1_81/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2602 vdd BUFX2_11/Y DFFPOSX1_79/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2603 DFFPOSX1_79/a_17_74# OAI22X1_14/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2604 DFFPOSX1_79/a_22_6# BUFX2_11/Y DFFPOSX1_79/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2605 DFFPOSX1_79/a_31_74# DFFPOSX1_79/a_2_6# DFFPOSX1_79/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2606 vdd DFFPOSX1_79/a_34_4# DFFPOSX1_79/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2607 DFFPOSX1_79/a_34_4# DFFPOSX1_79/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2608 DFFPOSX1_79/a_61_74# DFFPOSX1_79/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2609 DFFPOSX1_79/a_66_6# DFFPOSX1_79/a_2_6# DFFPOSX1_79/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2610 DFFPOSX1_79/a_76_84# BUFX2_11/Y DFFPOSX1_79/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2611 vdd out_MuxData[6] DFFPOSX1_79/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2612 gnd BUFX2_11/Y DFFPOSX1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2613 out_MuxData[6] DFFPOSX1_79/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2614 DFFPOSX1_79/a_17_6# OAI22X1_14/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2615 DFFPOSX1_79/a_22_6# DFFPOSX1_79/a_2_6# DFFPOSX1_79/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2616 DFFPOSX1_79/a_31_6# BUFX2_11/Y DFFPOSX1_79/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2617 gnd DFFPOSX1_79/a_34_4# DFFPOSX1_79/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2618 DFFPOSX1_79/a_34_4# DFFPOSX1_79/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2619 DFFPOSX1_79/a_61_6# DFFPOSX1_79/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2620 DFFPOSX1_79/a_66_6# BUFX2_11/Y DFFPOSX1_79/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2621 DFFPOSX1_79/a_76_6# DFFPOSX1_79/a_2_6# DFFPOSX1_79/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2622 gnd out_MuxData[6] DFFPOSX1_79/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2623 out_MuxData[6] DFFPOSX1_79/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2624 OAI22X1_13/a_9_54# INVX2_110/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2625 OAI22X1_13/Y INVX2_84/Y OAI22X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2626 OAI22X1_13/a_28_54# INVX2_99/Y OAI22X1_13/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2627 vdd XOR2X1_69/A OAI22X1_13/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2628 gnd INVX2_110/Y OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2629 OAI22X1_13/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2630 OAI22X1_13/Y INVX2_99/Y OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2631 OAI22X1_13/a_2_6# XOR2X1_69/A OAI22X1_13/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2632 INVX2_109/Y INVX2_109/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2633 INVX2_109/Y INVX2_109/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2634 vdd INVX2_61/Y DFFPOSX1_76/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2635 DFFPOSX1_76/a_17_74# OAI22X1_12/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2636 DFFPOSX1_76/a_22_6# INVX2_61/Y DFFPOSX1_76/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2637 DFFPOSX1_76/a_31_74# DFFPOSX1_76/a_2_6# DFFPOSX1_76/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2638 vdd DFFPOSX1_76/a_34_4# DFFPOSX1_76/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2639 DFFPOSX1_76/a_34_4# DFFPOSX1_76/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2640 DFFPOSX1_76/a_61_74# DFFPOSX1_76/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2641 DFFPOSX1_76/a_66_6# DFFPOSX1_76/a_2_6# DFFPOSX1_76/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2642 DFFPOSX1_76/a_76_84# INVX2_61/Y DFFPOSX1_76/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2643 vdd INVX2_109/A DFFPOSX1_76/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2644 gnd INVX2_61/Y DFFPOSX1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2645 INVX2_109/A DFFPOSX1_76/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2646 DFFPOSX1_76/a_17_6# OAI22X1_12/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2647 DFFPOSX1_76/a_22_6# DFFPOSX1_76/a_2_6# DFFPOSX1_76/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2648 DFFPOSX1_76/a_31_6# INVX2_61/Y DFFPOSX1_76/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2649 gnd DFFPOSX1_76/a_34_4# DFFPOSX1_76/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2650 DFFPOSX1_76/a_34_4# DFFPOSX1_76/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2651 DFFPOSX1_76/a_61_6# DFFPOSX1_76/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2652 DFFPOSX1_76/a_66_6# INVX2_61/Y DFFPOSX1_76/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2653 DFFPOSX1_76/a_76_6# DFFPOSX1_76/a_2_6# DFFPOSX1_76/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2654 gnd INVX2_109/A DFFPOSX1_76/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2655 INVX2_109/A DFFPOSX1_76/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2656 OAI22X1_12/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2657 OAI22X1_12/Y INVX2_109/Y OAI22X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2658 OAI22X1_12/a_28_54# INVX2_105/Y OAI22X1_12/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2659 vdd INVX2_62/Y OAI22X1_12/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2660 gnd BUFX2_4/Y OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2661 OAI22X1_12/a_2_6# INVX2_109/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2662 OAI22X1_12/Y INVX2_105/Y OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2663 OAI22X1_12/a_2_6# INVX2_62/Y OAI22X1_12/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2664 vdd INVX2_61/Y DFFPOSX1_75/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2665 DFFPOSX1_75/a_17_74# INVX2_107/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2666 DFFPOSX1_75/a_22_6# INVX2_61/Y DFFPOSX1_75/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2667 DFFPOSX1_75/a_31_74# DFFPOSX1_75/a_2_6# DFFPOSX1_75/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2668 vdd DFFPOSX1_75/a_34_4# DFFPOSX1_75/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2669 DFFPOSX1_75/a_34_4# DFFPOSX1_75/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2670 DFFPOSX1_75/a_61_74# DFFPOSX1_75/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2671 DFFPOSX1_75/a_66_6# DFFPOSX1_75/a_2_6# DFFPOSX1_75/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2672 DFFPOSX1_75/a_76_84# INVX2_61/Y DFFPOSX1_75/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2673 vdd AOI22X1_80/B DFFPOSX1_75/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2674 gnd INVX2_61/Y DFFPOSX1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2675 AOI22X1_80/B DFFPOSX1_75/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2676 DFFPOSX1_75/a_17_6# INVX2_107/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2677 DFFPOSX1_75/a_22_6# DFFPOSX1_75/a_2_6# DFFPOSX1_75/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2678 DFFPOSX1_75/a_31_6# INVX2_61/Y DFFPOSX1_75/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2679 gnd DFFPOSX1_75/a_34_4# DFFPOSX1_75/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2680 DFFPOSX1_75/a_34_4# DFFPOSX1_75/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2681 DFFPOSX1_75/a_61_6# DFFPOSX1_75/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2682 DFFPOSX1_75/a_66_6# INVX2_61/Y DFFPOSX1_75/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2683 DFFPOSX1_75/a_76_6# DFFPOSX1_75/a_2_6# DFFPOSX1_75/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2684 gnd AOI22X1_80/B DFFPOSX1_75/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2685 AOI22X1_80/B DFFPOSX1_75/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2686 INVX2_107/Y INVX2_107/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2687 INVX2_107/Y INVX2_107/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2688 NOR2X1_38/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2689 NOR2X1_38/Y INVX2_106/Y NOR2X1_38/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2690 NOR2X1_38/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2691 gnd INVX2_106/Y NOR2X1_38/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2692 vdd INVX2_62/Y AOI22X1_80/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2693 AOI22X1_80/a_2_54# AOI22X1_80/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2694 INVX2_107/A out_MemBData[5] AOI22X1_80/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2695 AOI22X1_80/a_2_54# BUFX2_8/Y INVX2_107/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2696 AOI22X1_80/a_11_6# INVX2_62/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2697 INVX2_107/A AOI22X1_80/B AOI22X1_80/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2698 AOI22X1_80/a_28_6# out_MemBData[5] INVX2_107/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2699 gnd BUFX2_8/Y AOI22X1_80/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2700 INVX2_106/Y INVX2_106/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2701 INVX2_106/Y INVX2_106/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2702 INVX2_105/Y out_MemBData[9] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2703 INVX2_105/Y out_MemBData[9] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2704 OAI21X1_70/a_9_54# NOR2X1_32/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2705 OAI21X1_69/C AND2X2_19/Y OAI21X1_70/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2706 vdd out_MemBData[9] OAI21X1_69/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2707 gnd NOR2X1_32/Y OAI21X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2708 OAI21X1_70/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2709 OAI21X1_69/C out_MemBData[9] OAI21X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2710 vdd BUFX2_10/Y DFFPOSX1_74/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2711 DFFPOSX1_74/a_17_74# OAI21X1_69/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2712 DFFPOSX1_74/a_22_6# BUFX2_10/Y DFFPOSX1_74/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2713 DFFPOSX1_74/a_31_74# DFFPOSX1_74/a_2_6# DFFPOSX1_74/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2714 vdd DFFPOSX1_74/a_34_4# DFFPOSX1_74/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2715 DFFPOSX1_74/a_34_4# DFFPOSX1_74/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2716 DFFPOSX1_74/a_61_74# DFFPOSX1_74/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2717 DFFPOSX1_74/a_66_6# DFFPOSX1_74/a_2_6# DFFPOSX1_74/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2718 DFFPOSX1_74/a_76_84# BUFX2_10/Y DFFPOSX1_74/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2719 vdd out_MemBData[9] DFFPOSX1_74/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2720 gnd BUFX2_10/Y DFFPOSX1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2721 out_MemBData[9] DFFPOSX1_74/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2722 DFFPOSX1_74/a_17_6# OAI21X1_69/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2723 DFFPOSX1_74/a_22_6# DFFPOSX1_74/a_2_6# DFFPOSX1_74/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2724 DFFPOSX1_74/a_31_6# BUFX2_10/Y DFFPOSX1_74/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2725 gnd DFFPOSX1_74/a_34_4# DFFPOSX1_74/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2726 DFFPOSX1_74/a_34_4# DFFPOSX1_74/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2727 DFFPOSX1_74/a_61_6# DFFPOSX1_74/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2728 DFFPOSX1_74/a_66_6# BUFX2_10/Y DFFPOSX1_74/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2729 DFFPOSX1_74/a_76_6# DFFPOSX1_74/a_2_6# DFFPOSX1_74/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2730 gnd out_MemBData[9] DFFPOSX1_74/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2731 out_MemBData[9] DFFPOSX1_74/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2732 OAI21X1_69/a_9_54# INVX2_93/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2733 OAI21X1_69/Y OR2X2_0/Y OAI21X1_69/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M2734 vdd OAI21X1_69/C OAI21X1_69/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2735 gnd INVX2_93/A OAI21X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M2736 OAI21X1_69/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2737 OAI21X1_69/Y OAI21X1_69/C OAI21X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2738 INVX2_93/A NOR2X1_36/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2739 vdd NOR2X1_30/Y INVX2_93/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2740 NAND2X1_33/a_9_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2741 INVX2_93/A NOR2X1_30/Y NAND2X1_33/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2742 INVX2_106/A NOR2X1_36/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2743 vdd NOR2X1_21/Y INVX2_106/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2744 NAND2X1_32/a_9_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2745 INVX2_106/A NOR2X1_21/Y NAND2X1_32/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2746 NOR2X1_34/a_9_54# con_count[3] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2747 NOR2X1_34/Y con_count[2] NOR2X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2748 NOR2X1_34/Y con_count[3] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2749 gnd con_count[2] NOR2X1_34/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2750 AND2X2_30/a_2_6# con_count[1] vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2751 vdd con_count[0] AND2X2_30/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2752 AND2X2_30/Y AND2X2_30/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2753 AND2X2_30/a_9_6# con_count[1] AND2X2_30/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M2754 gnd con_count[0] AND2X2_30/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2755 AND2X2_30/Y AND2X2_30/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2756 vdd con_count[1] HAX1_8/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M2757 HAX1_8/a_2_74# con_count[0] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2758 vdd HAX1_8/a_2_74# HAX1_10/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2759 HAX1_8/a_41_74# HAX1_8/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M2760 HAX1_8/a_49_54# con_count[0] HAX1_8/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2761 vdd con_count[1] HAX1_8/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2762 HAX1_8/YS HAX1_8/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2763 HAX1_8/a_9_6# con_count[1] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2764 HAX1_8/a_2_74# con_count[0] HAX1_8/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2765 gnd HAX1_8/a_2_74# HAX1_10/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M2766 HAX1_8/a_38_6# HAX1_8/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M2767 HAX1_8/a_41_74# con_count[0] HAX1_8/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2768 HAX1_8/a_38_6# con_count[1] HAX1_8/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2769 HAX1_8/YS HAX1_8/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2770 AND2X2_29/a_2_6# HAX1_8/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2771 vdd INVX2_72/Y AND2X2_29/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2772 AND2X2_29/Y AND2X2_29/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2773 AND2X2_29/a_9_6# HAX1_8/YS AND2X2_29/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M2774 gnd INVX2_72/Y AND2X2_29/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2775 AND2X2_29/Y AND2X2_29/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2776 INVX2_70/A NOR2X1_40/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M2777 vdd NAND3X1_29/Y INVX2_70/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2778 INVX2_70/A NOR2X1_33/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2779 NAND3X1_28/a_9_6# NOR2X1_40/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2780 NAND3X1_28/a_14_6# NAND3X1_29/Y NAND3X1_28/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M2781 INVX2_70/A NOR2X1_33/Y NAND3X1_28/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M2782 NOR2X1_33/a_9_54# con_count[6] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2783 NOR2X1_33/Y OR2X1_2/Y NOR2X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2784 NOR2X1_33/Y con_count[6] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M2785 gnd OR2X1_2/Y NOR2X1_33/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2786 vdd INVX2_43/Y DFFPOSX1_72/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2787 DFFPOSX1_72/a_17_74# INVX2_102/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2788 DFFPOSX1_72/a_22_6# INVX2_43/Y DFFPOSX1_72/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2789 DFFPOSX1_72/a_31_74# DFFPOSX1_72/a_2_6# DFFPOSX1_72/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2790 vdd DFFPOSX1_72/a_34_4# DFFPOSX1_72/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2791 DFFPOSX1_72/a_34_4# DFFPOSX1_72/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2792 DFFPOSX1_72/a_61_74# DFFPOSX1_72/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2793 DFFPOSX1_72/a_66_6# DFFPOSX1_72/a_2_6# DFFPOSX1_72/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2794 DFFPOSX1_72/a_76_84# INVX2_43/Y DFFPOSX1_72/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2795 vdd con_count[6] DFFPOSX1_72/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2796 gnd INVX2_43/Y DFFPOSX1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2797 con_count[6] DFFPOSX1_72/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2798 DFFPOSX1_72/a_17_6# INVX2_102/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2799 DFFPOSX1_72/a_22_6# DFFPOSX1_72/a_2_6# DFFPOSX1_72/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2800 DFFPOSX1_72/a_31_6# INVX2_43/Y DFFPOSX1_72/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2801 gnd DFFPOSX1_72/a_34_4# DFFPOSX1_72/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2802 DFFPOSX1_72/a_34_4# DFFPOSX1_72/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2803 DFFPOSX1_72/a_61_6# DFFPOSX1_72/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2804 DFFPOSX1_72/a_66_6# INVX2_43/Y DFFPOSX1_72/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2805 DFFPOSX1_72/a_76_6# DFFPOSX1_72/a_2_6# DFFPOSX1_72/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2806 gnd con_count[6] DFFPOSX1_72/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2807 con_count[6] DFFPOSX1_72/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2808 INVX2_102/Y INVX2_102/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2809 INVX2_102/Y INVX2_102/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2810 vdd out_MuxData[10] XOR2X1_74/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2811 XOR2X1_74/a_18_54# XOR2X1_74/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2812 XOR2X1_74/Y out_MuxData[10] XOR2X1_74/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2813 XOR2X1_74/a_35_54# XOR2X1_74/a_2_6# XOR2X1_74/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2814 vdd XOR2X1_74/B XOR2X1_74/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2815 XOR2X1_74/a_13_43# XOR2X1_74/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2816 gnd out_MuxData[10] XOR2X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2817 XOR2X1_74/a_18_6# XOR2X1_74/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2818 XOR2X1_74/Y XOR2X1_74/a_2_6# XOR2X1_74/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2819 XOR2X1_74/a_35_6# out_MuxData[10] XOR2X1_74/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2820 gnd XOR2X1_74/B XOR2X1_74/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2821 XOR2X1_74/a_13_43# XOR2X1_74/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2822 vdd OAI22X1_6/C XOR2X1_73/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2823 XOR2X1_73/a_18_54# XOR2X1_73/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2824 XOR2X1_72/B OAI22X1_6/C XOR2X1_73/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2825 XOR2X1_73/a_35_54# XOR2X1_73/a_2_6# XOR2X1_72/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2826 vdd XOR2X1_81/A XOR2X1_73/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2827 XOR2X1_73/a_13_43# XOR2X1_81/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2828 gnd OAI22X1_6/C XOR2X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2829 XOR2X1_73/a_18_6# XOR2X1_73/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2830 XOR2X1_72/B XOR2X1_73/a_2_6# XOR2X1_73/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2831 XOR2X1_73/a_35_6# OAI22X1_6/C XOR2X1_72/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2832 gnd XOR2X1_81/A XOR2X1_73/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2833 XOR2X1_73/a_13_43# XOR2X1_81/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2834 OAI22X1_6/C out_MuxData[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2835 OAI22X1_6/C out_MuxData[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2836 vdd out_MuxData[3] AOI22X1_76/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2837 AOI22X1_76/a_2_54# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2838 OAI21X1_89/A out_MuxData[9] AOI22X1_76/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2839 AOI22X1_76/a_2_54# XOR2X1_71/Y OAI21X1_89/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2840 AOI22X1_76/a_11_6# out_MuxData[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2841 OAI21X1_89/A out_MuxData[5] AOI22X1_76/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2842 AOI22X1_76/a_28_6# out_MuxData[9] OAI21X1_89/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2843 gnd XOR2X1_71/Y AOI22X1_76/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2844 vdd out_MuxData[5] XOR2X1_71/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2845 XOR2X1_71/a_18_54# XOR2X1_71/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2846 XOR2X1_71/Y out_MuxData[5] XOR2X1_71/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2847 XOR2X1_71/a_35_54# XOR2X1_71/a_2_6# XOR2X1_71/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2848 vdd INVX2_86/A XOR2X1_71/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2849 XOR2X1_71/a_13_43# INVX2_86/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2850 gnd out_MuxData[5] XOR2X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2851 XOR2X1_71/a_18_6# XOR2X1_71/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2852 XOR2X1_71/Y XOR2X1_71/a_2_6# XOR2X1_71/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2853 XOR2X1_71/a_35_6# out_MuxData[5] XOR2X1_71/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2854 gnd INVX2_86/A XOR2X1_71/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2855 XOR2X1_71/a_13_43# INVX2_86/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2856 out_MuxData[3] INVX2_86/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2857 out_MuxData[3] INVX2_86/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2858 vdd INVX2_86/Y XNOR2X1_46/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2859 XNOR2X1_46/a_18_54# XNOR2X1_46/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2860 XOR2X1_87/B XNOR2X1_46/a_2_6# XNOR2X1_46/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2861 XNOR2X1_46/a_35_54# INVX2_86/Y XOR2X1_87/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2862 vdd XOR2X1_70/Y XNOR2X1_46/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2863 XNOR2X1_46/a_12_41# XOR2X1_70/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2864 gnd INVX2_86/Y XNOR2X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2865 XNOR2X1_46/a_18_6# XNOR2X1_46/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2866 XOR2X1_87/B INVX2_86/Y XNOR2X1_46/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2867 XNOR2X1_46/a_35_6# XNOR2X1_46/a_2_6# XOR2X1_87/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2868 gnd XOR2X1_70/Y XNOR2X1_46/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2869 XNOR2X1_46/a_12_41# XOR2X1_70/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2870 vdd XOR2X1_70/Y AOI22X1_74/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2871 AOI22X1_74/a_2_54# out_MuxData[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2872 NOR2X1_42/A out_MuxData[0] AOI22X1_74/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2873 AOI22X1_74/a_2_54# XOR2X1_70/B NOR2X1_42/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2874 AOI22X1_74/a_11_6# XOR2X1_70/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2875 NOR2X1_42/A out_MuxData[3] AOI22X1_74/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2876 AOI22X1_74/a_28_6# out_MuxData[0] NOR2X1_42/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2877 gnd XOR2X1_70/B AOI22X1_74/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2878 vdd out_MuxData[0] XOR2X1_70/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2879 XOR2X1_70/a_18_54# XOR2X1_70/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2880 XOR2X1_70/Y out_MuxData[0] XOR2X1_70/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2881 XOR2X1_70/a_35_54# XOR2X1_70/a_2_6# XOR2X1_70/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2882 vdd XOR2X1_70/B XOR2X1_70/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2883 XOR2X1_70/a_13_43# XOR2X1_70/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2884 gnd out_MuxData[0] XOR2X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2885 XOR2X1_70/a_18_6# XOR2X1_70/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2886 XOR2X1_70/Y XOR2X1_70/a_2_6# XOR2X1_70/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2887 XOR2X1_70/a_35_6# out_MuxData[0] XOR2X1_70/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2888 gnd XOR2X1_70/B XOR2X1_70/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2889 XOR2X1_70/a_13_43# XOR2X1_70/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2890 vdd XOR2X1_69/A XOR2X1_69/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2891 XOR2X1_69/a_18_54# XOR2X1_69/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2892 XOR2X1_68/B XOR2X1_69/A XOR2X1_69/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2893 XOR2X1_69/a_35_54# XOR2X1_69/a_2_6# XOR2X1_68/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2894 vdd XOR2X1_69/B XOR2X1_69/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2895 XOR2X1_69/a_13_43# XOR2X1_69/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2896 gnd XOR2X1_69/A XOR2X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2897 XOR2X1_69/a_18_6# XOR2X1_69/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2898 XOR2X1_68/B XOR2X1_69/a_2_6# XOR2X1_69/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2899 XOR2X1_69/a_35_6# XOR2X1_69/A XOR2X1_68/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2900 gnd XOR2X1_69/B XOR2X1_69/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2901 XOR2X1_69/a_13_43# XOR2X1_69/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2902 vdd out_MuxData[5] XOR2X1_68/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2903 XOR2X1_68/a_18_54# XOR2X1_68/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2904 XOR2X1_67/B out_MuxData[5] XOR2X1_68/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M2905 XOR2X1_68/a_35_54# XOR2X1_68/a_2_6# XOR2X1_67/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2906 vdd XOR2X1_68/B XOR2X1_68/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2907 XOR2X1_68/a_13_43# XOR2X1_68/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2908 gnd out_MuxData[5] XOR2X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2909 XOR2X1_68/a_18_6# XOR2X1_68/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2910 XOR2X1_67/B XOR2X1_68/a_2_6# XOR2X1_68/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2911 XOR2X1_68/a_35_6# out_MuxData[5] XOR2X1_67/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2912 gnd XOR2X1_68/B XOR2X1_68/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2913 XOR2X1_68/a_13_43# XOR2X1_68/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2914 vdd BUFX2_10/Y DFFPOSX1_71/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2915 DFFPOSX1_71/a_17_74# OAI22X1_10/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2916 DFFPOSX1_71/a_22_6# BUFX2_10/Y DFFPOSX1_71/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2917 DFFPOSX1_71/a_31_74# DFFPOSX1_71/a_2_6# DFFPOSX1_71/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2918 vdd DFFPOSX1_71/a_34_4# DFFPOSX1_71/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2919 DFFPOSX1_71/a_34_4# DFFPOSX1_71/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2920 DFFPOSX1_71/a_61_74# DFFPOSX1_71/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2921 DFFPOSX1_71/a_66_6# DFFPOSX1_71/a_2_6# DFFPOSX1_71/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2922 DFFPOSX1_71/a_76_84# BUFX2_10/Y DFFPOSX1_71/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2923 vdd out_MuxData[9] DFFPOSX1_71/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2924 gnd BUFX2_10/Y DFFPOSX1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2925 out_MuxData[9] DFFPOSX1_71/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2926 DFFPOSX1_71/a_17_6# OAI22X1_10/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2927 DFFPOSX1_71/a_22_6# DFFPOSX1_71/a_2_6# DFFPOSX1_71/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2928 DFFPOSX1_71/a_31_6# BUFX2_10/Y DFFPOSX1_71/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2929 gnd DFFPOSX1_71/a_34_4# DFFPOSX1_71/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2930 DFFPOSX1_71/a_34_4# DFFPOSX1_71/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2931 DFFPOSX1_71/a_61_6# DFFPOSX1_71/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2932 DFFPOSX1_71/a_66_6# BUFX2_10/Y DFFPOSX1_71/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2933 DFFPOSX1_71/a_76_6# DFFPOSX1_71/a_2_6# DFFPOSX1_71/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2934 gnd out_MuxData[9] DFFPOSX1_71/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2935 out_MuxData[9] DFFPOSX1_71/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2936 OAI22X1_10/a_9_54# INVX2_109/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2937 OAI22X1_10/Y INVX2_84/Y OAI22X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M2938 OAI22X1_10/a_28_54# INVX2_99/Y OAI22X1_10/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M2939 vdd XOR2X1_69/B OAI22X1_10/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2940 gnd INVX2_109/Y OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M2941 OAI22X1_10/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2942 OAI22X1_10/Y INVX2_99/Y OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2943 OAI22X1_10/a_2_6# XOR2X1_69/B OAI22X1_10/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2944 vdd BUFX2_10/Y DFFPOSX1_70/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2945 DFFPOSX1_70/a_17_74# OAI22X1_13/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2946 DFFPOSX1_70/a_22_6# BUFX2_10/Y DFFPOSX1_70/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2947 DFFPOSX1_70/a_31_74# DFFPOSX1_70/a_2_6# DFFPOSX1_70/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2948 vdd DFFPOSX1_70/a_34_4# DFFPOSX1_70/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2949 DFFPOSX1_70/a_34_4# DFFPOSX1_70/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2950 DFFPOSX1_70/a_61_74# DFFPOSX1_70/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2951 DFFPOSX1_70/a_66_6# DFFPOSX1_70/a_2_6# DFFPOSX1_70/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2952 DFFPOSX1_70/a_76_84# BUFX2_10/Y DFFPOSX1_70/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2953 vdd out_MuxData[10] DFFPOSX1_70/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2954 gnd BUFX2_10/Y DFFPOSX1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2955 out_MuxData[10] DFFPOSX1_70/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2956 DFFPOSX1_70/a_17_6# OAI22X1_13/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2957 DFFPOSX1_70/a_22_6# DFFPOSX1_70/a_2_6# DFFPOSX1_70/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2958 DFFPOSX1_70/a_31_6# BUFX2_10/Y DFFPOSX1_70/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2959 gnd DFFPOSX1_70/a_34_4# DFFPOSX1_70/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2960 DFFPOSX1_70/a_34_4# DFFPOSX1_70/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2961 DFFPOSX1_70/a_61_6# DFFPOSX1_70/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2962 DFFPOSX1_70/a_66_6# BUFX2_10/Y DFFPOSX1_70/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M2963 DFFPOSX1_70/a_76_6# DFFPOSX1_70/a_2_6# DFFPOSX1_70/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2964 gnd out_MuxData[10] DFFPOSX1_70/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2965 out_MuxData[10] DFFPOSX1_70/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2966 vdd AOI22X1_80/B AOI22X1_72/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2967 AOI22X1_72/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2968 INVX2_98/A INVX2_99/A AOI22X1_72/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2969 AOI22X1_72/a_2_54# out_MuxData[5] INVX2_98/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2970 AOI22X1_72/a_11_6# AOI22X1_80/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2971 INVX2_98/A con_writeout AOI22X1_72/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2972 AOI22X1_72/a_28_6# INVX2_99/A INVX2_98/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2973 gnd out_MuxData[5] AOI22X1_72/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2974 vdd AOI22X1_69/B AOI22X1_70/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M2975 AOI22X1_70/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2976 INVX2_97/A INVX2_99/A AOI22X1_70/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M2977 AOI22X1_70/a_2_54# out_MuxData[4] INVX2_97/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2978 AOI22X1_70/a_11_6# AOI22X1_69/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2979 INVX2_97/A con_writeout AOI22X1_70/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M2980 AOI22X1_70/a_28_6# INVX2_99/A INVX2_97/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2981 gnd out_MuxData[4] AOI22X1_70/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2982 vdd INVX2_61/Y DFFPOSX1_68/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M2983 DFFPOSX1_68/a_17_74# INVX2_95/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2984 DFFPOSX1_68/a_22_6# INVX2_61/Y DFFPOSX1_68/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M2985 DFFPOSX1_68/a_31_74# DFFPOSX1_68/a_2_6# DFFPOSX1_68/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M2986 vdd DFFPOSX1_68/a_34_4# DFFPOSX1_68/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2987 DFFPOSX1_68/a_34_4# DFFPOSX1_68/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M2988 DFFPOSX1_68/a_61_74# DFFPOSX1_68/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M2989 DFFPOSX1_68/a_66_6# DFFPOSX1_68/a_2_6# DFFPOSX1_68/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M2990 DFFPOSX1_68/a_76_84# INVX2_61/Y DFFPOSX1_68/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2991 vdd AOI22X1_69/B DFFPOSX1_68/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2992 gnd INVX2_61/Y DFFPOSX1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M2993 AOI22X1_69/B DFFPOSX1_68/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M2994 DFFPOSX1_68/a_17_6# INVX2_95/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2995 DFFPOSX1_68/a_22_6# DFFPOSX1_68/a_2_6# DFFPOSX1_68/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2996 DFFPOSX1_68/a_31_6# INVX2_61/Y DFFPOSX1_68/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M2997 gnd DFFPOSX1_68/a_34_4# DFFPOSX1_68/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2998 DFFPOSX1_68/a_34_4# DFFPOSX1_68/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M2999 DFFPOSX1_68/a_61_6# DFFPOSX1_68/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3000 DFFPOSX1_68/a_66_6# INVX2_61/Y DFFPOSX1_68/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3001 DFFPOSX1_68/a_76_6# DFFPOSX1_68/a_2_6# DFFPOSX1_68/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3002 gnd AOI22X1_69/B DFFPOSX1_68/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3003 AOI22X1_69/B DFFPOSX1_68/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3004 vdd INVX2_62/Y AOI22X1_69/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3005 AOI22X1_69/a_2_54# AOI22X1_69/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3006 INVX2_95/A out_MemBData[4] AOI22X1_69/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3007 AOI22X1_69/a_2_54# BUFX2_8/Y INVX2_95/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3008 AOI22X1_69/a_11_6# INVX2_62/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3009 INVX2_95/A AOI22X1_69/B AOI22X1_69/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3010 AOI22X1_69/a_28_6# out_MemBData[4] INVX2_95/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3011 gnd BUFX2_8/Y AOI22X1_69/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3012 vdd BUFX2_10/Y DFFPOSX1_67/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3013 DFFPOSX1_67/a_17_74# OAI21X1_65/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3014 DFFPOSX1_67/a_22_6# BUFX2_10/Y DFFPOSX1_67/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3015 DFFPOSX1_67/a_31_74# DFFPOSX1_67/a_2_6# DFFPOSX1_67/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3016 vdd DFFPOSX1_67/a_34_4# DFFPOSX1_67/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3017 DFFPOSX1_67/a_34_4# DFFPOSX1_67/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3018 DFFPOSX1_67/a_61_74# DFFPOSX1_67/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3019 DFFPOSX1_67/a_66_6# DFFPOSX1_67/a_2_6# DFFPOSX1_67/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3020 DFFPOSX1_67/a_76_84# BUFX2_10/Y DFFPOSX1_67/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3021 vdd out_MemBData[12] DFFPOSX1_67/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3022 gnd BUFX2_10/Y DFFPOSX1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3023 out_MemBData[12] DFFPOSX1_67/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3024 DFFPOSX1_67/a_17_6# OAI21X1_65/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3025 DFFPOSX1_67/a_22_6# DFFPOSX1_67/a_2_6# DFFPOSX1_67/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3026 DFFPOSX1_67/a_31_6# BUFX2_10/Y DFFPOSX1_67/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3027 gnd DFFPOSX1_67/a_34_4# DFFPOSX1_67/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3028 DFFPOSX1_67/a_34_4# DFFPOSX1_67/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3029 DFFPOSX1_67/a_61_6# DFFPOSX1_67/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3030 DFFPOSX1_67/a_66_6# BUFX2_10/Y DFFPOSX1_67/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3031 DFFPOSX1_67/a_76_6# DFFPOSX1_67/a_2_6# DFFPOSX1_67/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3032 gnd out_MemBData[12] DFFPOSX1_67/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3033 out_MemBData[12] DFFPOSX1_67/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3034 OAI21X1_66/a_9_54# NOR2X1_23/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3035 OAI21X1_65/C AND2X2_19/Y OAI21X1_66/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3036 vdd out_MemBData[12] OAI21X1_65/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3037 gnd NOR2X1_23/Y OAI21X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3038 OAI21X1_66/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3039 OAI21X1_65/C out_MemBData[12] OAI21X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3040 OAI21X1_65/a_9_54# INVX2_92/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3041 OAI21X1_65/Y OR2X2_0/Y OAI21X1_65/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3042 vdd OAI21X1_65/C OAI21X1_65/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3043 gnd INVX2_92/A OAI21X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3044 OAI21X1_65/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3045 OAI21X1_65/Y OAI21X1_65/C OAI21X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3046 INVX2_92/A NOR2X1_35/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3047 vdd NOR2X1_31/Y INVX2_92/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3048 NAND2X1_30/a_9_6# NOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3049 INVX2_92/A NOR2X1_31/Y NAND2X1_30/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3050 NOR2X1_31/a_9_54# con_count[1] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3051 NOR2X1_31/Y con_count[0] NOR2X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3052 NOR2X1_31/Y con_count[1] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3053 gnd con_count[0] NOR2X1_31/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3054 vdd INVX2_43/Y DFFPOSX1_66/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3055 DFFPOSX1_66/a_17_74# INVX2_89/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3056 DFFPOSX1_66/a_22_6# INVX2_43/Y DFFPOSX1_66/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3057 DFFPOSX1_66/a_31_74# DFFPOSX1_66/a_2_6# DFFPOSX1_66/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3058 vdd DFFPOSX1_66/a_34_4# DFFPOSX1_66/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3059 DFFPOSX1_66/a_34_4# DFFPOSX1_66/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3060 DFFPOSX1_66/a_61_74# DFFPOSX1_66/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3061 DFFPOSX1_66/a_66_6# DFFPOSX1_66/a_2_6# DFFPOSX1_66/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3062 DFFPOSX1_66/a_76_84# INVX2_43/Y DFFPOSX1_66/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3063 vdd con_count[1] DFFPOSX1_66/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3064 gnd INVX2_43/Y DFFPOSX1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3065 con_count[1] DFFPOSX1_66/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3066 DFFPOSX1_66/a_17_6# INVX2_89/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3067 DFFPOSX1_66/a_22_6# DFFPOSX1_66/a_2_6# DFFPOSX1_66/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3068 DFFPOSX1_66/a_31_6# INVX2_43/Y DFFPOSX1_66/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3069 gnd DFFPOSX1_66/a_34_4# DFFPOSX1_66/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3070 DFFPOSX1_66/a_34_4# DFFPOSX1_66/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3071 DFFPOSX1_66/a_61_6# DFFPOSX1_66/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3072 DFFPOSX1_66/a_66_6# INVX2_43/Y DFFPOSX1_66/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3073 DFFPOSX1_66/a_76_6# DFFPOSX1_66/a_2_6# DFFPOSX1_66/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3074 gnd con_count[1] DFFPOSX1_66/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3075 con_count[1] DFFPOSX1_66/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3076 vdd BUFX2_9/Y DFFPOSX1_65/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3077 DFFPOSX1_65/a_17_74# AND2X2_29/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3078 DFFPOSX1_65/a_22_6# BUFX2_9/Y DFFPOSX1_65/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3079 DFFPOSX1_65/a_31_74# DFFPOSX1_65/a_2_6# DFFPOSX1_65/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3080 vdd DFFPOSX1_65/a_34_4# DFFPOSX1_65/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3081 DFFPOSX1_65/a_34_4# DFFPOSX1_65/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3082 DFFPOSX1_65/a_61_74# DFFPOSX1_65/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3083 DFFPOSX1_65/a_66_6# DFFPOSX1_65/a_2_6# DFFPOSX1_65/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3084 DFFPOSX1_65/a_76_84# BUFX2_9/Y DFFPOSX1_65/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3085 vdd AOI22X1_68/C DFFPOSX1_65/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3086 gnd BUFX2_9/Y DFFPOSX1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3087 AOI22X1_68/C DFFPOSX1_65/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3088 DFFPOSX1_65/a_17_6# AND2X2_29/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3089 DFFPOSX1_65/a_22_6# DFFPOSX1_65/a_2_6# DFFPOSX1_65/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3090 DFFPOSX1_65/a_31_6# BUFX2_9/Y DFFPOSX1_65/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3091 gnd DFFPOSX1_65/a_34_4# DFFPOSX1_65/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3092 DFFPOSX1_65/a_34_4# DFFPOSX1_65/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3093 DFFPOSX1_65/a_61_6# DFFPOSX1_65/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3094 DFFPOSX1_65/a_66_6# BUFX2_9/Y DFFPOSX1_65/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3095 DFFPOSX1_65/a_76_6# DFFPOSX1_65/a_2_6# DFFPOSX1_65/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3096 gnd AOI22X1_68/C DFFPOSX1_65/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3097 AOI22X1_68/C DFFPOSX1_65/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3098 AND2X2_27/a_2_6# HAX1_7/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3099 vdd INVX2_72/Y AND2X2_27/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3100 AND2X2_27/Y AND2X2_27/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3101 AND2X2_27/a_9_6# HAX1_7/YS AND2X2_27/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M3102 gnd INVX2_72/Y AND2X2_27/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3103 AND2X2_27/Y AND2X2_27/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3104 vdd BUFX2_9/Y DFFPOSX1_64/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3105 DFFPOSX1_64/a_17_74# AND2X2_27/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3106 DFFPOSX1_64/a_22_6# BUFX2_9/Y DFFPOSX1_64/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3107 DFFPOSX1_64/a_31_74# DFFPOSX1_64/a_2_6# DFFPOSX1_64/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3108 vdd DFFPOSX1_64/a_34_4# DFFPOSX1_64/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3109 DFFPOSX1_64/a_34_4# DFFPOSX1_64/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3110 DFFPOSX1_64/a_61_74# DFFPOSX1_64/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3111 DFFPOSX1_64/a_66_6# DFFPOSX1_64/a_2_6# DFFPOSX1_64/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3112 DFFPOSX1_64/a_76_84# BUFX2_9/Y DFFPOSX1_64/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3113 vdd AOI22X1_67/C DFFPOSX1_64/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3114 gnd BUFX2_9/Y DFFPOSX1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3115 AOI22X1_67/C DFFPOSX1_64/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3116 DFFPOSX1_64/a_17_6# AND2X2_27/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3117 DFFPOSX1_64/a_22_6# DFFPOSX1_64/a_2_6# DFFPOSX1_64/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3118 DFFPOSX1_64/a_31_6# BUFX2_9/Y DFFPOSX1_64/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3119 gnd DFFPOSX1_64/a_34_4# DFFPOSX1_64/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3120 DFFPOSX1_64/a_34_4# DFFPOSX1_64/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3121 DFFPOSX1_64/a_61_6# DFFPOSX1_64/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3122 DFFPOSX1_64/a_66_6# BUFX2_9/Y DFFPOSX1_64/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3123 DFFPOSX1_64/a_76_6# DFFPOSX1_64/a_2_6# DFFPOSX1_64/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3124 gnd AOI22X1_67/C DFFPOSX1_64/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3125 AOI22X1_67/C DFFPOSX1_64/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3126 vdd XOR2X1_74/Y AOI22X1_78/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3127 AOI22X1_78/a_2_54# out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3128 NOR2X1_29/A out_MuxData[10] AOI22X1_78/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3129 AOI22X1_78/a_2_54# XOR2X1_74/B NOR2X1_29/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3130 AOI22X1_78/a_11_6# XOR2X1_74/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3131 NOR2X1_29/A out_MuxData[9] AOI22X1_78/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3132 AOI22X1_78/a_28_6# out_MuxData[10] NOR2X1_29/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3133 gnd XOR2X1_74/B AOI22X1_78/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3134 vdd out_MuxData[0] AOI22X1_77/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3135 AOI22X1_77/a_2_54# out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3136 NOR2X1_29/B out_MuxData[12] AOI22X1_77/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3137 AOI22X1_77/a_2_54# XOR2X1_72/B NOR2X1_29/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3138 AOI22X1_77/a_11_6# out_MuxData[0] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3139 NOR2X1_29/B out_MuxData[1] AOI22X1_77/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3140 AOI22X1_77/a_28_6# out_MuxData[12] NOR2X1_29/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3141 gnd XOR2X1_72/B AOI22X1_77/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3142 vdd out_MuxData[12] XOR2X1_72/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3143 XOR2X1_72/a_18_54# XOR2X1_72/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3144 XOR2X1_74/B out_MuxData[12] XOR2X1_72/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3145 XOR2X1_72/a_35_54# XOR2X1_72/a_2_6# XOR2X1_74/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3146 vdd XOR2X1_72/B XOR2X1_72/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3147 XOR2X1_72/a_13_43# XOR2X1_72/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3148 gnd out_MuxData[12] XOR2X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3149 XOR2X1_72/a_18_6# XOR2X1_72/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3150 XOR2X1_74/B XOR2X1_72/a_2_6# XOR2X1_72/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3151 XOR2X1_72/a_35_6# out_MuxData[12] XOR2X1_74/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3152 gnd XOR2X1_72/B XOR2X1_72/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3153 XOR2X1_72/a_13_43# XOR2X1_72/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3154 vdd out_MuxData[10] AOI22X1_75/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3155 AOI22X1_75/a_2_54# out_MuxData[12] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3156 OAI21X1_68/A out_MuxData[0] AOI22X1_75/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3157 AOI22X1_75/a_2_54# XOR2X1_66/Y OAI21X1_68/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3158 AOI22X1_75/a_11_6# out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3159 OAI21X1_68/A out_MuxData[12] AOI22X1_75/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3160 AOI22X1_75/a_28_6# out_MuxData[0] OAI21X1_68/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3161 gnd XOR2X1_66/Y AOI22X1_75/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3162 NAND3X1_27/B OAI21X1_68/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3163 vdd OAI21X1_68/B NAND3X1_27/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3164 NAND2X1_31/a_9_6# OAI21X1_68/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3165 NAND3X1_27/B OAI21X1_68/B NAND2X1_31/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3166 OAI21X1_68/a_9_54# OAI21X1_68/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3167 XNOR2X1_45/A OAI21X1_68/B OAI21X1_68/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3168 vdd NAND3X1_27/B XNOR2X1_45/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3169 gnd OAI21X1_68/A OAI21X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3170 OAI21X1_68/a_2_6# OAI21X1_68/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3171 XNOR2X1_45/A NAND3X1_27/B OAI21X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3172 NAND3X1_27/Y AND2X2_28/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M3173 vdd NAND3X1_27/B NAND3X1_27/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3174 NAND3X1_27/Y AND2X2_28/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3175 NAND3X1_27/a_9_6# AND2X2_28/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M3176 NAND3X1_27/a_14_6# NAND3X1_27/B NAND3X1_27/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M3177 NAND3X1_27/Y AND2X2_28/B NAND3X1_27/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M3178 AND2X2_28/a_2_6# AND2X2_28/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3179 vdd AND2X2_28/B AND2X2_28/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3180 AND2X2_28/Y AND2X2_28/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3181 AND2X2_28/a_9_6# AND2X2_28/A AND2X2_28/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M3182 gnd AND2X2_28/B AND2X2_28/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3183 AND2X2_28/Y AND2X2_28/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3184 vdd XNOR2X1_45/A XNOR2X1_45/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3185 XNOR2X1_45/a_18_54# XNOR2X1_45/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3186 XNOR2X1_45/Y XNOR2X1_45/a_2_6# XNOR2X1_45/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3187 XNOR2X1_45/a_35_54# XNOR2X1_45/A XNOR2X1_45/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3188 vdd AND2X2_28/Y XNOR2X1_45/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3189 XNOR2X1_45/a_12_41# AND2X2_28/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3190 gnd XNOR2X1_45/A XNOR2X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3191 XNOR2X1_45/a_18_6# XNOR2X1_45/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3192 XNOR2X1_45/Y XNOR2X1_45/A XNOR2X1_45/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3193 XNOR2X1_45/a_35_6# XNOR2X1_45/a_2_6# XNOR2X1_45/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3194 gnd AND2X2_28/Y XNOR2X1_45/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3195 XNOR2X1_45/a_12_41# AND2X2_28/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3196 vdd XOR2X1_69/A XNOR2X1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3197 XNOR2X1_44/a_18_54# XNOR2X1_44/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3198 XOR2X1_55/B XNOR2X1_44/a_2_6# XNOR2X1_44/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3199 XNOR2X1_44/a_35_54# XOR2X1_69/A XOR2X1_55/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3200 vdd XOR2X1_62/Y XNOR2X1_44/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3201 XNOR2X1_44/a_12_41# XOR2X1_62/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3202 gnd XOR2X1_69/A XNOR2X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3203 XNOR2X1_44/a_18_6# XNOR2X1_44/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3204 XOR2X1_55/B XOR2X1_69/A XNOR2X1_44/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3205 XNOR2X1_44/a_35_6# XNOR2X1_44/a_2_6# XOR2X1_55/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3206 gnd XOR2X1_62/Y XNOR2X1_44/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3207 XNOR2X1_44/a_12_41# XOR2X1_62/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3208 vdd XOR2X1_67/B AOI22X1_73/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3209 AOI22X1_73/a_2_54# out_MuxData[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3210 AOI21X1_7/B out_MuxData[2] AOI22X1_73/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3211 AOI22X1_73/a_2_54# XOR2X1_67/Y AOI21X1_7/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3212 AOI22X1_73/a_11_6# XOR2X1_67/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3213 AOI21X1_7/B out_MuxData[3] AOI22X1_73/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3214 AOI22X1_73/a_28_6# out_MuxData[2] AOI21X1_7/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3215 gnd XOR2X1_67/Y AOI22X1_73/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3216 vdd INVX2_86/A XOR2X1_67/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3217 XOR2X1_67/a_18_54# XOR2X1_67/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3218 XOR2X1_67/Y INVX2_86/A XOR2X1_67/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3219 XOR2X1_67/a_35_54# XOR2X1_67/a_2_6# XOR2X1_67/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3220 vdd XOR2X1_67/B XOR2X1_67/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3221 XOR2X1_67/a_13_43# XOR2X1_67/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3222 gnd INVX2_86/A XOR2X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3223 XOR2X1_67/a_18_6# XOR2X1_67/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3224 XOR2X1_67/Y XOR2X1_67/a_2_6# XOR2X1_67/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3225 XOR2X1_67/a_35_6# INVX2_86/A XOR2X1_67/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3226 gnd XOR2X1_67/B XOR2X1_67/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3227 XOR2X1_67/a_13_43# XOR2X1_67/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3228 vdd INVX2_85/Y XNOR2X1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3229 XNOR2X1_43/a_18_54# XNOR2X1_43/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3230 AND2X2_36/A XNOR2X1_43/a_2_6# XNOR2X1_43/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3231 XNOR2X1_43/a_35_54# INVX2_85/Y AND2X2_36/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3232 vdd XOR2X1_67/Y XNOR2X1_43/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3233 XNOR2X1_43/a_12_41# XOR2X1_67/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3234 gnd INVX2_85/Y XNOR2X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3235 XNOR2X1_43/a_18_6# XNOR2X1_43/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3236 AND2X2_36/A INVX2_85/Y XNOR2X1_43/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3237 XNOR2X1_43/a_35_6# XNOR2X1_43/a_2_6# AND2X2_36/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3238 gnd XOR2X1_67/Y XNOR2X1_43/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3239 XNOR2X1_43/a_12_41# XOR2X1_67/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3240 INVX2_99/Y INVX2_99/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3241 INVX2_99/Y INVX2_99/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3242 vdd BUFX2_11/Y DFFPOSX1_69/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3243 DFFPOSX1_69/a_17_74# INVX2_97/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3244 DFFPOSX1_69/a_22_6# BUFX2_11/Y DFFPOSX1_69/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3245 DFFPOSX1_69/a_31_74# DFFPOSX1_69/a_2_6# DFFPOSX1_69/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3246 vdd DFFPOSX1_69/a_34_4# DFFPOSX1_69/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3247 DFFPOSX1_69/a_34_4# DFFPOSX1_69/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3248 DFFPOSX1_69/a_61_74# DFFPOSX1_69/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3249 DFFPOSX1_69/a_66_6# DFFPOSX1_69/a_2_6# DFFPOSX1_69/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3250 DFFPOSX1_69/a_76_84# BUFX2_11/Y DFFPOSX1_69/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3251 vdd out_MuxData[4] DFFPOSX1_69/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3252 gnd BUFX2_11/Y DFFPOSX1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3253 out_MuxData[4] DFFPOSX1_69/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3254 DFFPOSX1_69/a_17_6# INVX2_97/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3255 DFFPOSX1_69/a_22_6# DFFPOSX1_69/a_2_6# DFFPOSX1_69/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3256 DFFPOSX1_69/a_31_6# BUFX2_11/Y DFFPOSX1_69/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3257 gnd DFFPOSX1_69/a_34_4# DFFPOSX1_69/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3258 DFFPOSX1_69/a_34_4# DFFPOSX1_69/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3259 DFFPOSX1_69/a_61_6# DFFPOSX1_69/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3260 DFFPOSX1_69/a_66_6# BUFX2_11/Y DFFPOSX1_69/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3261 DFFPOSX1_69/a_76_6# DFFPOSX1_69/a_2_6# DFFPOSX1_69/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3262 gnd out_MuxData[4] DFFPOSX1_69/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3263 out_MuxData[4] DFFPOSX1_69/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3264 INVX2_98/Y INVX2_98/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3265 INVX2_98/Y INVX2_98/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3266 vdd AOI22X1_62/B AOI22X1_71/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3267 AOI22X1_71/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3268 INVX2_82/A INVX2_99/A AOI22X1_71/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3269 AOI22X1_71/a_2_54# out_MuxData[12] INVX2_82/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3270 AOI22X1_71/a_11_6# AOI22X1_62/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3271 INVX2_82/A con_writeout AOI22X1_71/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3272 AOI22X1_71/a_28_6# INVX2_99/A INVX2_82/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3273 gnd out_MuxData[12] AOI22X1_71/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3274 INVX2_97/Y INVX2_97/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3275 INVX2_97/Y INVX2_97/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3276 INVX2_96/Y INVX2_96/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3277 INVX2_96/Y INVX2_96/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3278 INVX2_95/Y INVX2_95/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3279 INVX2_95/Y INVX2_95/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3280 NOR2X1_32/a_9_54# INVX2_62/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3281 NOR2X1_32/Y INVX2_93/Y NOR2X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3282 NOR2X1_32/Y INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3283 gnd INVX2_93/Y NOR2X1_32/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3284 INVX2_94/Y INVX2_94/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3285 INVX2_94/Y INVX2_94/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3286 INVX2_93/Y INVX2_93/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3287 INVX2_93/Y INVX2_93/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3288 OAI21X1_67/a_9_54# INVX2_94/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3289 OAI21X1_67/Y OR2X2_0/Y OAI21X1_67/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3290 vdd OAI21X1_67/C OAI21X1_67/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3291 gnd INVX2_94/A OAI21X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3292 OAI21X1_67/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3293 OAI21X1_67/Y OAI21X1_67/C OAI21X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3294 INVX2_92/Y INVX2_92/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3295 INVX2_92/Y INVX2_92/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3296 vdd in_clka BUFX2_11/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3297 BUFX2_11/Y BUFX2_11/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3298 gnd in_clka BUFX2_11/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M3299 BUFX2_11/Y BUFX2_11/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3300 INVX2_94/A NOR2X1_35/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3301 vdd NOR2X1_30/Y INVX2_94/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3302 NAND2X1_29/a_9_6# NOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3303 INVX2_94/A NOR2X1_30/Y NAND2X1_29/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3304 NOR2X1_30/a_9_54# INVX2_91/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3305 NOR2X1_30/Y con_count[1] NOR2X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3306 NOR2X1_30/Y INVX2_91/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3307 gnd con_count[1] NOR2X1_30/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3308 INVX2_91/Y con_count[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3309 INVX2_91/Y con_count[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3310 INVX2_90/Y con_count[1] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3311 INVX2_90/Y con_count[1] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3312 INVX2_89/Y INVX2_89/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3313 INVX2_89/Y INVX2_89/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3314 vdd con_count[1] AOI22X1_68/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3315 AOI22X1_68/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3316 INVX2_89/A INVX2_126/A AOI22X1_68/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3317 AOI22X1_68/a_2_54# AOI22X1_68/C INVX2_89/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3318 AOI22X1_68/a_11_6# con_count[1] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3319 INVX2_89/A INVX2_126/Y AOI22X1_68/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3320 AOI22X1_68/a_28_6# INVX2_126/A INVX2_89/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3321 gnd AOI22X1_68/C AOI22X1_68/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3322 vdd con_count[7] HAX1_7/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M3323 HAX1_7/a_2_74# HAX1_7/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3324 vdd HAX1_7/a_2_74# HAX1_7/YC vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3325 HAX1_7/a_41_74# HAX1_7/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M3326 HAX1_7/a_49_54# HAX1_7/B HAX1_7/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3327 vdd con_count[7] HAX1_7/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3328 HAX1_7/YS HAX1_7/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3329 HAX1_7/a_9_6# con_count[7] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3330 HAX1_7/a_2_74# HAX1_7/B HAX1_7/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3331 gnd HAX1_7/a_2_74# HAX1_7/YC Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M3332 HAX1_7/a_38_6# HAX1_7/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M3333 HAX1_7/a_41_74# HAX1_7/B HAX1_7/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3334 HAX1_7/a_38_6# con_count[7] HAX1_7/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3335 HAX1_7/YS HAX1_7/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3336 OR2X1_2/a_9_54# con_count[8] OR2X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M3337 vdd con_count[7] OR2X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3338 OR2X1_2/Y OR2X1_2/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3339 OR2X1_2/a_2_54# con_count[8] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3340 gnd con_count[7] OR2X1_2/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3341 OR2X1_2/Y OR2X1_2/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3342 vdd con_count[7] AOI22X1_67/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3343 AOI22X1_67/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3344 INVX2_88/A INVX2_126/A AOI22X1_67/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3345 AOI22X1_67/a_2_54# AOI22X1_67/C INVX2_88/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3346 AOI22X1_67/a_11_6# con_count[7] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3347 INVX2_88/A INVX2_126/Y AOI22X1_67/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3348 AOI22X1_67/a_28_6# INVX2_126/A INVX2_88/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3349 gnd AOI22X1_67/C AOI22X1_67/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3350 INVX2_88/Y INVX2_88/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3351 INVX2_88/Y INVX2_88/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3352 vdd XOR2X1_69/B XNOR2X1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3353 XNOR2X1_42/a_18_54# XNOR2X1_42/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3354 XOR2X1_58/B XNOR2X1_42/a_2_6# XNOR2X1_42/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3355 XNOR2X1_42/a_35_54# XOR2X1_69/B XOR2X1_58/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3356 vdd XOR2X1_74/Y XNOR2X1_42/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3357 XNOR2X1_42/a_12_41# XOR2X1_74/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3358 gnd XOR2X1_69/B XNOR2X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3359 XNOR2X1_42/a_18_6# XNOR2X1_42/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3360 XOR2X1_58/B XOR2X1_69/B XNOR2X1_42/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3361 XNOR2X1_42/a_35_6# XNOR2X1_42/a_2_6# XOR2X1_58/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3362 gnd XOR2X1_74/Y XNOR2X1_42/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3363 XNOR2X1_42/a_12_41# XOR2X1_74/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3364 vdd NOR2X1_29/B XNOR2X1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3365 XNOR2X1_41/a_18_54# XNOR2X1_41/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3366 XNOR2X1_41/Y XNOR2X1_41/a_2_6# XNOR2X1_41/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3367 XNOR2X1_41/a_35_54# NOR2X1_29/B XNOR2X1_41/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3368 vdd NOR2X1_29/A XNOR2X1_41/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3369 XNOR2X1_41/a_12_41# NOR2X1_29/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3370 gnd NOR2X1_29/B XNOR2X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3371 XNOR2X1_41/a_18_6# XNOR2X1_41/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3372 XNOR2X1_41/Y NOR2X1_29/B XNOR2X1_41/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3373 XNOR2X1_41/a_35_6# XNOR2X1_41/a_2_6# XNOR2X1_41/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3374 gnd NOR2X1_29/A XNOR2X1_41/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3375 XNOR2X1_41/a_12_41# NOR2X1_29/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3376 NOR2X1_29/a_9_54# NOR2X1_29/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3377 XOR2X1_65/B NOR2X1_29/B NOR2X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3378 XOR2X1_65/B NOR2X1_29/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3379 gnd NOR2X1_29/B XOR2X1_65/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3380 vdd out_MuxData[12] XOR2X1_66/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3381 XOR2X1_66/a_18_54# XOR2X1_66/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3382 XOR2X1_66/Y out_MuxData[12] XOR2X1_66/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3383 XOR2X1_66/a_35_54# XOR2X1_66/a_2_6# XOR2X1_66/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3384 vdd out_MuxData[10] XOR2X1_66/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3385 XOR2X1_66/a_13_43# out_MuxData[10] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3386 gnd out_MuxData[12] XOR2X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3387 XOR2X1_66/a_18_6# XOR2X1_66/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3388 XOR2X1_66/Y XOR2X1_66/a_2_6# XOR2X1_66/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3389 XOR2X1_66/a_35_6# out_MuxData[12] XOR2X1_66/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3390 gnd out_MuxData[10] XOR2X1_66/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3391 XOR2X1_66/a_13_43# out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3392 vdd OAI22X1_6/C XNOR2X1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3393 XNOR2X1_40/a_18_54# XNOR2X1_40/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3394 AND2X2_28/B XNOR2X1_40/a_2_6# XNOR2X1_40/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3395 XNOR2X1_40/a_35_54# OAI22X1_6/C AND2X2_28/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3396 vdd XOR2X1_66/Y XNOR2X1_40/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3397 XNOR2X1_40/a_12_41# XOR2X1_66/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3398 gnd OAI22X1_6/C XNOR2X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3399 XNOR2X1_40/a_18_6# XNOR2X1_40/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3400 AND2X2_28/B OAI22X1_6/C XNOR2X1_40/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3401 XNOR2X1_40/a_35_6# XNOR2X1_40/a_2_6# AND2X2_28/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3402 gnd XOR2X1_66/Y XNOR2X1_40/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3403 XNOR2X1_40/a_12_41# XOR2X1_66/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3404 vdd NOR2X1_28/B XNOR2X1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3405 XNOR2X1_39/a_18_54# XNOR2X1_39/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3406 OAI21X1_68/B XNOR2X1_39/a_2_6# XNOR2X1_39/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3407 XNOR2X1_39/a_35_54# NOR2X1_28/B OAI21X1_68/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3408 vdd NOR2X1_28/A XNOR2X1_39/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3409 XNOR2X1_39/a_12_41# NOR2X1_28/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3410 gnd NOR2X1_28/B XNOR2X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3411 XNOR2X1_39/a_18_6# XNOR2X1_39/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3412 OAI21X1_68/B NOR2X1_28/B XNOR2X1_39/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3413 XNOR2X1_39/a_35_6# XNOR2X1_39/a_2_6# OAI21X1_68/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3414 gnd NOR2X1_28/A XNOR2X1_39/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3415 XNOR2X1_39/a_12_41# NOR2X1_28/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3416 OAI21X1_64/a_9_54# OAI21X1_68/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3417 XOR2X1_57/A OAI21X1_68/B OAI21X1_64/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3418 vdd NAND3X1_27/Y XOR2X1_57/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3419 gnd OAI21X1_68/A OAI21X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3420 OAI21X1_64/a_2_6# OAI21X1_68/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3421 XOR2X1_57/A NAND3X1_27/Y OAI21X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3422 vdd AND2X2_28/B XOR2X1_63/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3423 XOR2X1_63/a_18_54# XOR2X1_63/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3424 XOR2X1_63/Y AND2X2_28/B XOR2X1_63/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3425 XOR2X1_63/a_35_54# XOR2X1_63/a_2_6# XOR2X1_63/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3426 vdd AND2X2_28/A XOR2X1_63/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3427 XOR2X1_63/a_13_43# AND2X2_28/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3428 gnd AND2X2_28/B XOR2X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3429 XOR2X1_63/a_18_6# XOR2X1_63/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3430 XOR2X1_63/Y XOR2X1_63/a_2_6# XOR2X1_63/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3431 XOR2X1_63/a_35_6# AND2X2_28/B XOR2X1_63/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3432 gnd AND2X2_28/A XOR2X1_63/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3433 XOR2X1_63/a_13_43# AND2X2_28/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3434 INVX2_87/Y out_MuxData[11] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3435 INVX2_87/Y out_MuxData[11] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3436 INVX2_86/Y INVX2_86/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3437 INVX2_86/Y INVX2_86/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3438 vdd out_MuxData[11] XOR2X1_62/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3439 XOR2X1_62/a_18_54# XOR2X1_62/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3440 XOR2X1_62/Y out_MuxData[11] XOR2X1_62/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3441 XOR2X1_62/a_35_54# XOR2X1_62/a_2_6# XOR2X1_62/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3442 vdd XOR2X1_62/B XOR2X1_62/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3443 XOR2X1_62/a_13_43# XOR2X1_62/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3444 gnd out_MuxData[11] XOR2X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3445 XOR2X1_62/a_18_6# XOR2X1_62/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3446 XOR2X1_62/Y XOR2X1_62/a_2_6# XOR2X1_62/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3447 XOR2X1_62/a_35_6# out_MuxData[11] XOR2X1_62/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3448 gnd XOR2X1_62/B XOR2X1_62/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3449 XOR2X1_62/a_13_43# XOR2X1_62/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3450 vdd XOR2X1_62/B AOI22X1_64/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3451 AOI22X1_64/a_2_54# out_MuxData[11] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3452 AOI21X1_6/B out_MuxData[10] AOI22X1_64/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3453 AOI22X1_64/a_2_54# XOR2X1_62/Y AOI21X1_6/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3454 AOI22X1_64/a_11_6# XOR2X1_62/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3455 AOI21X1_6/B out_MuxData[11] AOI22X1_64/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3456 AOI22X1_64/a_28_6# out_MuxData[10] AOI21X1_6/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3457 gnd XOR2X1_62/Y AOI22X1_64/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3458 INVX2_85/Y out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3459 INVX2_85/Y out_MuxData[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3460 vdd BUFX2_11/Y DFFPOSX1_63/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3461 DFFPOSX1_63/a_17_74# INVX2_98/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3462 DFFPOSX1_63/a_22_6# BUFX2_11/Y DFFPOSX1_63/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3463 DFFPOSX1_63/a_31_74# DFFPOSX1_63/a_2_6# DFFPOSX1_63/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3464 vdd DFFPOSX1_63/a_34_4# DFFPOSX1_63/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3465 DFFPOSX1_63/a_34_4# DFFPOSX1_63/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3466 DFFPOSX1_63/a_61_74# DFFPOSX1_63/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3467 DFFPOSX1_63/a_66_6# DFFPOSX1_63/a_2_6# DFFPOSX1_63/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3468 DFFPOSX1_63/a_76_84# BUFX2_11/Y DFFPOSX1_63/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3469 vdd out_MuxData[5] DFFPOSX1_63/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3470 gnd BUFX2_11/Y DFFPOSX1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3471 out_MuxData[5] DFFPOSX1_63/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3472 DFFPOSX1_63/a_17_6# INVX2_98/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3473 DFFPOSX1_63/a_22_6# DFFPOSX1_63/a_2_6# DFFPOSX1_63/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3474 DFFPOSX1_63/a_31_6# BUFX2_11/Y DFFPOSX1_63/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3475 gnd DFFPOSX1_63/a_34_4# DFFPOSX1_63/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3476 DFFPOSX1_63/a_34_4# DFFPOSX1_63/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3477 DFFPOSX1_63/a_61_6# DFFPOSX1_63/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3478 DFFPOSX1_63/a_66_6# BUFX2_11/Y DFFPOSX1_63/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3479 DFFPOSX1_63/a_76_6# DFFPOSX1_63/a_2_6# DFFPOSX1_63/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3480 gnd out_MuxData[5] DFFPOSX1_63/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3481 out_MuxData[5] DFFPOSX1_63/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3482 vdd BUFX2_10/Y DFFPOSX1_62/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3483 DFFPOSX1_62/a_17_74# INVX2_83/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3484 DFFPOSX1_62/a_22_6# BUFX2_10/Y DFFPOSX1_62/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3485 DFFPOSX1_62/a_31_74# DFFPOSX1_62/a_2_6# DFFPOSX1_62/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3486 vdd DFFPOSX1_62/a_34_4# DFFPOSX1_62/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3487 DFFPOSX1_62/a_34_4# DFFPOSX1_62/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3488 DFFPOSX1_62/a_61_74# DFFPOSX1_62/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3489 DFFPOSX1_62/a_66_6# DFFPOSX1_62/a_2_6# DFFPOSX1_62/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3490 DFFPOSX1_62/a_76_84# BUFX2_10/Y DFFPOSX1_62/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3491 vdd out_MuxData[13] DFFPOSX1_62/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3492 gnd BUFX2_10/Y DFFPOSX1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3493 out_MuxData[13] DFFPOSX1_62/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3494 DFFPOSX1_62/a_17_6# INVX2_83/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3495 DFFPOSX1_62/a_22_6# DFFPOSX1_62/a_2_6# DFFPOSX1_62/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3496 DFFPOSX1_62/a_31_6# BUFX2_10/Y DFFPOSX1_62/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3497 gnd DFFPOSX1_62/a_34_4# DFFPOSX1_62/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3498 DFFPOSX1_62/a_34_4# DFFPOSX1_62/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3499 DFFPOSX1_62/a_61_6# DFFPOSX1_62/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3500 DFFPOSX1_62/a_66_6# BUFX2_10/Y DFFPOSX1_62/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3501 DFFPOSX1_62/a_76_6# DFFPOSX1_62/a_2_6# DFFPOSX1_62/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3502 gnd out_MuxData[13] DFFPOSX1_62/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3503 out_MuxData[13] DFFPOSX1_62/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3504 vdd BUFX2_10/Y DFFPOSX1_61/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3505 DFFPOSX1_61/a_17_74# INVX2_82/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3506 DFFPOSX1_61/a_22_6# BUFX2_10/Y DFFPOSX1_61/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3507 DFFPOSX1_61/a_31_74# DFFPOSX1_61/a_2_6# DFFPOSX1_61/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3508 vdd DFFPOSX1_61/a_34_4# DFFPOSX1_61/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3509 DFFPOSX1_61/a_34_4# DFFPOSX1_61/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3510 DFFPOSX1_61/a_61_74# DFFPOSX1_61/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3511 DFFPOSX1_61/a_66_6# DFFPOSX1_61/a_2_6# DFFPOSX1_61/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3512 DFFPOSX1_61/a_76_84# BUFX2_10/Y DFFPOSX1_61/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3513 vdd out_MuxData[12] DFFPOSX1_61/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3514 gnd BUFX2_10/Y DFFPOSX1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3515 out_MuxData[12] DFFPOSX1_61/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3516 DFFPOSX1_61/a_17_6# INVX2_82/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3517 DFFPOSX1_61/a_22_6# DFFPOSX1_61/a_2_6# DFFPOSX1_61/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3518 DFFPOSX1_61/a_31_6# BUFX2_10/Y DFFPOSX1_61/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3519 gnd DFFPOSX1_61/a_34_4# DFFPOSX1_61/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3520 DFFPOSX1_61/a_34_4# DFFPOSX1_61/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3521 DFFPOSX1_61/a_61_6# DFFPOSX1_61/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3522 DFFPOSX1_61/a_66_6# BUFX2_10/Y DFFPOSX1_61/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3523 DFFPOSX1_61/a_76_6# DFFPOSX1_61/a_2_6# DFFPOSX1_61/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3524 gnd out_MuxData[12] DFFPOSX1_61/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3525 out_MuxData[12] DFFPOSX1_61/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3526 INVX2_82/Y INVX2_82/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3527 INVX2_82/Y INVX2_82/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3528 vdd INVX2_61/Y DFFPOSX1_60/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3529 DFFPOSX1_60/a_17_74# INVX2_96/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3530 DFFPOSX1_60/a_22_6# INVX2_61/Y DFFPOSX1_60/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3531 DFFPOSX1_60/a_31_74# DFFPOSX1_60/a_2_6# DFFPOSX1_60/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3532 vdd DFFPOSX1_60/a_34_4# DFFPOSX1_60/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3533 DFFPOSX1_60/a_34_4# DFFPOSX1_60/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3534 DFFPOSX1_60/a_61_74# DFFPOSX1_60/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3535 DFFPOSX1_60/a_66_6# DFFPOSX1_60/a_2_6# DFFPOSX1_60/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3536 DFFPOSX1_60/a_76_84# INVX2_61/Y DFFPOSX1_60/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3537 vdd AOI22X1_62/B DFFPOSX1_60/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3538 gnd INVX2_61/Y DFFPOSX1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3539 AOI22X1_62/B DFFPOSX1_60/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3540 DFFPOSX1_60/a_17_6# INVX2_96/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3541 DFFPOSX1_60/a_22_6# DFFPOSX1_60/a_2_6# DFFPOSX1_60/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3542 DFFPOSX1_60/a_31_6# INVX2_61/Y DFFPOSX1_60/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3543 gnd DFFPOSX1_60/a_34_4# DFFPOSX1_60/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3544 DFFPOSX1_60/a_34_4# DFFPOSX1_60/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3545 DFFPOSX1_60/a_61_6# DFFPOSX1_60/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3546 DFFPOSX1_60/a_66_6# INVX2_61/Y DFFPOSX1_60/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3547 DFFPOSX1_60/a_76_6# DFFPOSX1_60/a_2_6# DFFPOSX1_60/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3548 gnd AOI22X1_62/B DFFPOSX1_60/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3549 AOI22X1_62/B DFFPOSX1_60/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3550 vdd INVX2_62/Y AOI22X1_62/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3551 AOI22X1_62/a_2_54# AOI22X1_62/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3552 INVX2_96/A out_MemBData[12] AOI22X1_62/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3553 AOI22X1_62/a_2_54# BUFX2_8/Y INVX2_96/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3554 AOI22X1_62/a_11_6# INVX2_62/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3555 INVX2_96/A AOI22X1_62/B AOI22X1_62/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3556 AOI22X1_62/a_28_6# out_MemBData[12] INVX2_96/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3557 gnd BUFX2_8/Y AOI22X1_62/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3558 NOR2X1_25/a_9_54# INVX2_62/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3559 NOR2X1_25/Y INVX2_94/Y NOR2X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3560 NOR2X1_25/Y INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3561 gnd INVX2_94/Y NOR2X1_25/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3562 OAI21X1_63/a_9_54# NOR2X1_25/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3563 OAI21X1_67/C AND2X2_19/Y OAI21X1_63/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3564 vdd out_MemBData[13] OAI21X1_67/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3565 gnd NOR2X1_25/Y OAI21X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3566 OAI21X1_63/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3567 OAI21X1_67/C out_MemBData[13] OAI21X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3568 vdd BUFX2_10/Y DFFPOSX1_58/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3569 DFFPOSX1_58/a_17_74# OAI21X1_67/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3570 DFFPOSX1_58/a_22_6# BUFX2_10/Y DFFPOSX1_58/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3571 DFFPOSX1_58/a_31_74# DFFPOSX1_58/a_2_6# DFFPOSX1_58/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3572 vdd DFFPOSX1_58/a_34_4# DFFPOSX1_58/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3573 DFFPOSX1_58/a_34_4# DFFPOSX1_58/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3574 DFFPOSX1_58/a_61_74# DFFPOSX1_58/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3575 DFFPOSX1_58/a_66_6# DFFPOSX1_58/a_2_6# DFFPOSX1_58/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3576 DFFPOSX1_58/a_76_84# BUFX2_10/Y DFFPOSX1_58/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3577 vdd out_MemBData[13] DFFPOSX1_58/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3578 gnd BUFX2_10/Y DFFPOSX1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3579 out_MemBData[13] DFFPOSX1_58/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3580 DFFPOSX1_58/a_17_6# OAI21X1_67/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3581 DFFPOSX1_58/a_22_6# DFFPOSX1_58/a_2_6# DFFPOSX1_58/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3582 DFFPOSX1_58/a_31_6# BUFX2_10/Y DFFPOSX1_58/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3583 gnd DFFPOSX1_58/a_34_4# DFFPOSX1_58/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3584 DFFPOSX1_58/a_34_4# DFFPOSX1_58/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3585 DFFPOSX1_58/a_61_6# DFFPOSX1_58/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3586 DFFPOSX1_58/a_66_6# BUFX2_10/Y DFFPOSX1_58/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3587 DFFPOSX1_58/a_76_6# DFFPOSX1_58/a_2_6# DFFPOSX1_58/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3588 gnd out_MemBData[13] DFFPOSX1_58/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3589 out_MemBData[13] DFFPOSX1_58/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3590 vdd in_clka BUFX2_10/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3591 BUFX2_10/Y BUFX2_10/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3592 gnd in_clka BUFX2_10/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M3593 BUFX2_10/Y BUFX2_10/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3594 INVX2_25/A NOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3595 vdd NOR2X1_30/Y INVX2_25/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3596 NAND2X1_27/a_9_6# NOR2X1_34/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3597 INVX2_25/A NOR2X1_30/Y NAND2X1_27/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3598 INVX2_71/A NOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3599 vdd NOR2X1_31/Y INVX2_71/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3600 NAND2X1_24/a_9_6# NOR2X1_34/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3601 INVX2_71/A NOR2X1_31/Y NAND2X1_24/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3602 NOR2X1_22/a_9_54# INVX2_90/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3603 NOR2X1_22/Y INVX2_91/Y NOR2X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3604 NOR2X1_22/Y INVX2_90/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3605 gnd INVX2_91/Y NOR2X1_22/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3606 NOR2X1_21/a_9_54# INVX2_90/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3607 NOR2X1_21/Y con_count[0] NOR2X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3608 NOR2X1_21/Y INVX2_90/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3609 gnd con_count[0] NOR2X1_21/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3610 vdd in_clka BUFX2_9/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3611 BUFX2_9/Y BUFX2_9/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3612 gnd in_clka BUFX2_9/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M3613 BUFX2_9/Y BUFX2_9/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3614 AND2X2_26/a_2_6# INVX2_91/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3615 vdd INVX2_72/Y AND2X2_26/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3616 AND2X2_26/Y AND2X2_26/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3617 AND2X2_26/a_9_6# INVX2_91/Y AND2X2_26/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M3618 gnd INVX2_72/Y AND2X2_26/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3619 AND2X2_26/Y AND2X2_26/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3620 vdd BUFX2_9/Y DFFPOSX1_57/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3621 DFFPOSX1_57/a_17_74# AND2X2_26/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3622 DFFPOSX1_57/a_22_6# BUFX2_9/Y DFFPOSX1_57/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3623 DFFPOSX1_57/a_31_74# DFFPOSX1_57/a_2_6# DFFPOSX1_57/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3624 vdd DFFPOSX1_57/a_34_4# DFFPOSX1_57/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3625 DFFPOSX1_57/a_34_4# DFFPOSX1_57/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3626 DFFPOSX1_57/a_61_74# DFFPOSX1_57/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3627 DFFPOSX1_57/a_66_6# DFFPOSX1_57/a_2_6# DFFPOSX1_57/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3628 DFFPOSX1_57/a_76_84# BUFX2_9/Y DFFPOSX1_57/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3629 vdd AOI22X1_60/C DFFPOSX1_57/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3630 gnd BUFX2_9/Y DFFPOSX1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3631 AOI22X1_60/C DFFPOSX1_57/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3632 DFFPOSX1_57/a_17_6# AND2X2_26/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3633 DFFPOSX1_57/a_22_6# DFFPOSX1_57/a_2_6# DFFPOSX1_57/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3634 DFFPOSX1_57/a_31_6# BUFX2_9/Y DFFPOSX1_57/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3635 gnd DFFPOSX1_57/a_34_4# DFFPOSX1_57/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3636 DFFPOSX1_57/a_34_4# DFFPOSX1_57/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3637 DFFPOSX1_57/a_61_6# DFFPOSX1_57/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3638 DFFPOSX1_57/a_66_6# BUFX2_9/Y DFFPOSX1_57/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3639 DFFPOSX1_57/a_76_6# DFFPOSX1_57/a_2_6# DFFPOSX1_57/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3640 gnd AOI22X1_60/C DFFPOSX1_57/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3641 AOI22X1_60/C DFFPOSX1_57/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3642 AND2X2_25/a_2_6# XOR2X1_59/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3643 vdd INVX2_72/Y AND2X2_25/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3644 AND2X2_25/Y AND2X2_25/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3645 AND2X2_25/a_9_6# XOR2X1_59/Y AND2X2_25/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M3646 gnd INVX2_72/Y AND2X2_25/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3647 AND2X2_25/Y AND2X2_25/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3648 vdd HAX1_7/YC XOR2X1_59/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3649 XOR2X1_59/a_18_54# XOR2X1_59/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3650 XOR2X1_59/Y HAX1_7/YC XOR2X1_59/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3651 XOR2X1_59/a_35_54# XOR2X1_59/a_2_6# XOR2X1_59/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3652 vdd con_count[8] XOR2X1_59/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3653 XOR2X1_59/a_13_43# con_count[8] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3654 gnd HAX1_7/YC XOR2X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3655 XOR2X1_59/a_18_6# XOR2X1_59/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3656 XOR2X1_59/Y XOR2X1_59/a_2_6# XOR2X1_59/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3657 XOR2X1_59/a_35_6# HAX1_7/YC XOR2X1_59/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3658 gnd con_count[8] XOR2X1_59/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3659 XOR2X1_59/a_13_43# con_count[8] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3660 vdd BUFX2_9/Y DFFPOSX1_56/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3661 DFFPOSX1_56/a_17_74# AND2X2_25/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3662 DFFPOSX1_56/a_22_6# BUFX2_9/Y DFFPOSX1_56/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3663 DFFPOSX1_56/a_31_74# DFFPOSX1_56/a_2_6# DFFPOSX1_56/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3664 vdd DFFPOSX1_56/a_34_4# DFFPOSX1_56/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3665 DFFPOSX1_56/a_34_4# DFFPOSX1_56/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3666 DFFPOSX1_56/a_61_74# DFFPOSX1_56/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3667 DFFPOSX1_56/a_66_6# DFFPOSX1_56/a_2_6# DFFPOSX1_56/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3668 DFFPOSX1_56/a_76_84# BUFX2_9/Y DFFPOSX1_56/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3669 vdd AOI22X1_59/C DFFPOSX1_56/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3670 gnd BUFX2_9/Y DFFPOSX1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3671 AOI22X1_59/C DFFPOSX1_56/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3672 DFFPOSX1_56/a_17_6# AND2X2_25/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3673 DFFPOSX1_56/a_22_6# DFFPOSX1_56/a_2_6# DFFPOSX1_56/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3674 DFFPOSX1_56/a_31_6# BUFX2_9/Y DFFPOSX1_56/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3675 gnd DFFPOSX1_56/a_34_4# DFFPOSX1_56/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3676 DFFPOSX1_56/a_34_4# DFFPOSX1_56/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3677 DFFPOSX1_56/a_61_6# DFFPOSX1_56/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3678 DFFPOSX1_56/a_66_6# BUFX2_9/Y DFFPOSX1_56/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3679 DFFPOSX1_56/a_76_6# DFFPOSX1_56/a_2_6# DFFPOSX1_56/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3680 gnd AOI22X1_59/C DFFPOSX1_56/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3681 AOI22X1_59/C DFFPOSX1_56/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3682 vdd INVX2_43/Y DFFPOSX1_55/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3683 DFFPOSX1_55/a_17_74# INVX2_88/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3684 DFFPOSX1_55/a_22_6# INVX2_43/Y DFFPOSX1_55/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3685 DFFPOSX1_55/a_31_74# DFFPOSX1_55/a_2_6# DFFPOSX1_55/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3686 vdd DFFPOSX1_55/a_34_4# DFFPOSX1_55/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3687 DFFPOSX1_55/a_34_4# DFFPOSX1_55/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3688 DFFPOSX1_55/a_61_74# DFFPOSX1_55/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3689 DFFPOSX1_55/a_66_6# DFFPOSX1_55/a_2_6# DFFPOSX1_55/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3690 DFFPOSX1_55/a_76_84# INVX2_43/Y DFFPOSX1_55/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3691 vdd con_count[7] DFFPOSX1_55/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3692 gnd INVX2_43/Y DFFPOSX1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3693 con_count[7] DFFPOSX1_55/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3694 DFFPOSX1_55/a_17_6# INVX2_88/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3695 DFFPOSX1_55/a_22_6# DFFPOSX1_55/a_2_6# DFFPOSX1_55/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3696 DFFPOSX1_55/a_31_6# INVX2_43/Y DFFPOSX1_55/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3697 gnd DFFPOSX1_55/a_34_4# DFFPOSX1_55/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3698 DFFPOSX1_55/a_34_4# DFFPOSX1_55/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3699 DFFPOSX1_55/a_61_6# DFFPOSX1_55/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3700 DFFPOSX1_55/a_66_6# INVX2_43/Y DFFPOSX1_55/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3701 DFFPOSX1_55/a_76_6# DFFPOSX1_55/a_2_6# DFFPOSX1_55/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3702 gnd con_count[7] DFFPOSX1_55/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3703 con_count[7] DFFPOSX1_55/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3704 NAND2X1_28/Y AOI22X1_58/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3705 vdd XNOR2X1_41/Y NAND2X1_28/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3706 NAND2X1_28/a_9_6# AOI22X1_58/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3707 NAND2X1_28/Y XNOR2X1_41/Y NAND2X1_28/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3708 vdd XOR2X1_65/A XOR2X1_65/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3709 XOR2X1_65/a_18_54# XOR2X1_65/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3710 XOR2X1_65/Y XOR2X1_65/A XOR2X1_65/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3711 XOR2X1_65/a_35_54# XOR2X1_65/a_2_6# XOR2X1_65/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3712 vdd XOR2X1_65/B XOR2X1_65/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3713 XOR2X1_65/a_13_43# XOR2X1_65/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3714 gnd XOR2X1_65/A XOR2X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3715 XOR2X1_65/a_18_6# XOR2X1_65/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3716 XOR2X1_65/Y XOR2X1_65/a_2_6# XOR2X1_65/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3717 XOR2X1_65/a_35_6# XOR2X1_65/A XOR2X1_65/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3718 gnd XOR2X1_65/B XOR2X1_65/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3719 XOR2X1_65/a_13_43# XOR2X1_65/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3720 vdd out_MuxData[8] XOR2X1_64/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3721 XOR2X1_64/a_18_54# XOR2X1_64/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3722 XOR2X1_64/Y out_MuxData[8] XOR2X1_64/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3723 XOR2X1_64/a_35_54# XOR2X1_64/a_2_6# XOR2X1_64/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3724 vdd XOR2X1_64/B XOR2X1_64/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3725 XOR2X1_64/a_13_43# XOR2X1_64/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3726 gnd out_MuxData[8] XOR2X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3727 XOR2X1_64/a_18_6# XOR2X1_64/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3728 XOR2X1_64/Y XOR2X1_64/a_2_6# XOR2X1_64/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3729 XOR2X1_64/a_35_6# out_MuxData[8] XOR2X1_64/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3730 gnd XOR2X1_64/B XOR2X1_64/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3731 XOR2X1_64/a_13_43# XOR2X1_64/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3732 vdd XOR2X1_64/B AOI22X1_66/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3733 AOI22X1_66/a_2_54# out_MuxData[8] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3734 NOR2X1_28/A out_MuxData[11] AOI22X1_66/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3735 AOI22X1_66/a_2_54# XOR2X1_64/Y NOR2X1_28/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3736 AOI22X1_66/a_11_6# XOR2X1_64/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3737 NOR2X1_28/A out_MuxData[8] AOI22X1_66/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3738 AOI22X1_66/a_28_6# out_MuxData[11] NOR2X1_28/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3739 gnd XOR2X1_64/Y AOI22X1_66/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3740 NOR2X1_28/a_9_54# NOR2X1_28/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3741 NOR2X1_28/Y NOR2X1_28/B NOR2X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3742 NOR2X1_28/Y NOR2X1_28/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3743 gnd NOR2X1_28/B NOR2X1_28/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3744 vdd INVX2_87/Y XNOR2X1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3745 XNOR2X1_38/a_18_54# XNOR2X1_38/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3746 AND2X2_28/A XNOR2X1_38/a_2_6# XNOR2X1_38/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3747 XNOR2X1_38/a_35_54# INVX2_87/Y AND2X2_28/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3748 vdd XOR2X1_64/Y XNOR2X1_38/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3749 XNOR2X1_38/a_12_41# XOR2X1_64/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3750 gnd INVX2_87/Y XNOR2X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3751 XNOR2X1_38/a_18_6# XNOR2X1_38/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3752 AND2X2_28/A INVX2_87/Y XNOR2X1_38/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3753 XNOR2X1_38/a_35_6# XNOR2X1_38/a_2_6# AND2X2_28/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3754 gnd XOR2X1_64/Y XNOR2X1_38/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3755 XNOR2X1_38/a_12_41# XOR2X1_64/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3756 vdd XOR2X1_65/Y AOI22X1_65/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3757 AOI22X1_65/a_2_54# INVX2_94/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3758 AND2X2_20/A INVX2_75/Y AOI22X1_65/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3759 AOI22X1_65/a_2_54# XOR2X1_61/Y AND2X2_20/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3760 AOI22X1_65/a_11_6# XOR2X1_65/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3761 AND2X2_20/A INVX2_94/Y AOI22X1_65/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3762 AOI22X1_65/a_28_6# INVX2_75/Y AND2X2_20/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3763 gnd XOR2X1_61/Y AOI22X1_65/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3764 vdd XOR2X1_61/A XOR2X1_61/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3765 XOR2X1_61/a_18_54# XOR2X1_61/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3766 XOR2X1_61/Y XOR2X1_61/A XOR2X1_61/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3767 XOR2X1_61/a_35_54# XOR2X1_61/a_2_6# XOR2X1_61/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3768 vdd NOR2X1_27/Y XOR2X1_61/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3769 XOR2X1_61/a_13_43# NOR2X1_27/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3770 gnd XOR2X1_61/A XOR2X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3771 XOR2X1_61/a_18_6# XOR2X1_61/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3772 XOR2X1_61/Y XOR2X1_61/a_2_6# XOR2X1_61/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3773 XOR2X1_61/a_35_6# XOR2X1_61/A XOR2X1_61/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3774 gnd NOR2X1_27/Y XOR2X1_61/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3775 XOR2X1_61/a_13_43# NOR2X1_27/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3776 NOR2X1_27/a_9_54# NOR2X1_27/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3777 NOR2X1_27/Y AOI21X1_6/B NOR2X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3778 NOR2X1_27/Y NOR2X1_27/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3779 gnd AOI21X1_6/B NOR2X1_27/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3780 vdd INVX2_50/Y XNOR2X1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3781 XNOR2X1_37/a_18_54# XNOR2X1_37/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3782 XOR2X1_62/B XNOR2X1_37/a_2_6# XNOR2X1_37/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3783 XNOR2X1_37/a_35_54# INVX2_50/Y XOR2X1_62/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3784 vdd XOR2X1_60/Y XNOR2X1_37/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3785 XNOR2X1_37/a_12_41# XOR2X1_60/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3786 gnd INVX2_50/Y XNOR2X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3787 XNOR2X1_37/a_18_6# XNOR2X1_37/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3788 XOR2X1_62/B INVX2_50/Y XNOR2X1_37/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3789 XNOR2X1_37/a_35_6# XNOR2X1_37/a_2_6# XOR2X1_62/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3790 gnd XOR2X1_60/Y XNOR2X1_37/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3791 XNOR2X1_37/a_12_41# XOR2X1_60/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3792 vdd XOR2X1_81/A XOR2X1_60/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3793 XOR2X1_60/a_18_54# XOR2X1_60/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3794 XOR2X1_60/Y XOR2X1_81/A XOR2X1_60/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3795 XOR2X1_60/a_35_54# XOR2X1_60/a_2_6# XOR2X1_60/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3796 vdd INVX2_85/Y XOR2X1_60/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3797 XOR2X1_60/a_13_43# INVX2_85/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3798 gnd XOR2X1_81/A XOR2X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3799 XOR2X1_60/a_18_6# XOR2X1_60/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3800 XOR2X1_60/Y XOR2X1_60/a_2_6# XOR2X1_60/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3801 XOR2X1_60/a_35_6# XOR2X1_81/A XOR2X1_60/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3802 gnd INVX2_85/Y XOR2X1_60/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3803 XOR2X1_60/a_13_43# INVX2_85/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3804 INVX2_84/Y con_writeout vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3805 INVX2_84/Y con_writeout gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3806 INVX2_83/Y INVX2_83/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3807 INVX2_83/Y INVX2_83/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3808 vdd AOI22X1_61/B AOI22X1_63/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3809 AOI22X1_63/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3810 INVX2_83/A INVX2_99/A AOI22X1_63/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3811 AOI22X1_63/a_2_54# out_MuxData[13] INVX2_83/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3812 AOI22X1_63/a_11_6# AOI22X1_61/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3813 INVX2_83/A con_writeout AOI22X1_63/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3814 AOI22X1_63/a_28_6# INVX2_99/A INVX2_83/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3815 gnd out_MuxData[13] AOI22X1_63/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3816 NOR2X1_26/a_9_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3817 INVX2_99/A INVX2_62/Y NOR2X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3818 INVX2_99/A con_writeout gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3819 gnd INVX2_62/Y INVX2_99/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3820 vdd INVX2_61/Y DFFPOSX1_59/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3821 DFFPOSX1_59/a_17_74# INVX2_81/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3822 DFFPOSX1_59/a_22_6# INVX2_61/Y DFFPOSX1_59/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3823 DFFPOSX1_59/a_31_74# DFFPOSX1_59/a_2_6# DFFPOSX1_59/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3824 vdd DFFPOSX1_59/a_34_4# DFFPOSX1_59/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3825 DFFPOSX1_59/a_34_4# DFFPOSX1_59/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3826 DFFPOSX1_59/a_61_74# DFFPOSX1_59/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3827 DFFPOSX1_59/a_66_6# DFFPOSX1_59/a_2_6# DFFPOSX1_59/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3828 DFFPOSX1_59/a_76_84# INVX2_61/Y DFFPOSX1_59/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3829 vdd AOI22X1_61/B DFFPOSX1_59/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3830 gnd INVX2_61/Y DFFPOSX1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3831 AOI22X1_61/B DFFPOSX1_59/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3832 DFFPOSX1_59/a_17_6# INVX2_81/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3833 DFFPOSX1_59/a_22_6# DFFPOSX1_59/a_2_6# DFFPOSX1_59/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3834 DFFPOSX1_59/a_31_6# INVX2_61/Y DFFPOSX1_59/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3835 gnd DFFPOSX1_59/a_34_4# DFFPOSX1_59/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3836 DFFPOSX1_59/a_34_4# DFFPOSX1_59/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3837 DFFPOSX1_59/a_61_6# DFFPOSX1_59/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3838 DFFPOSX1_59/a_66_6# INVX2_61/Y DFFPOSX1_59/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3839 DFFPOSX1_59/a_76_6# DFFPOSX1_59/a_2_6# DFFPOSX1_59/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3840 gnd AOI22X1_61/B DFFPOSX1_59/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3841 AOI22X1_61/B DFFPOSX1_59/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3842 INVX2_81/Y INVX2_81/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3843 INVX2_81/Y INVX2_81/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3844 vdd con_restart AOI22X1_61/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3845 AOI22X1_61/a_2_54# AOI22X1_61/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3846 INVX2_81/A out_MemBData[13] AOI22X1_61/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3847 AOI22X1_61/a_2_54# BUFX2_7/Y INVX2_81/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3848 AOI22X1_61/a_11_6# con_restart gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3849 INVX2_81/A AOI22X1_61/B AOI22X1_61/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3850 AOI22X1_61/a_28_6# out_MemBData[13] INVX2_81/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3851 gnd BUFX2_7/Y AOI22X1_61/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3852 NOR2X1_24/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3853 NOR2X1_24/Y INVX2_75/Y NOR2X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3854 NOR2X1_24/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3855 gnd INVX2_75/Y NOR2X1_24/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3856 OAI21X1_62/a_9_54# NOR2X1_24/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3857 OAI21X1_62/Y AND2X2_19/Y OAI21X1_62/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3858 vdd out_MemBData[14] OAI21X1_62/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3859 gnd NOR2X1_24/Y OAI21X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3860 OAI21X1_62/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3861 OAI21X1_62/Y out_MemBData[14] OAI21X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3862 OAI21X1_61/a_9_54# INVX2_75/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3863 OAI21X1_61/Y OR2X2_0/Y OAI21X1_61/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3864 vdd OAI21X1_62/Y OAI21X1_61/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3865 gnd INVX2_75/A OAI21X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3866 OAI21X1_61/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3867 OAI21X1_61/Y OAI21X1_62/Y OAI21X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3868 NOR2X1_23/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3869 NOR2X1_23/Y INVX2_92/Y NOR2X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3870 NOR2X1_23/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M3871 gnd INVX2_92/Y NOR2X1_23/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3872 INVX2_26/A NOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3873 vdd NOR2X1_22/Y INVX2_26/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3874 NAND2X1_26/a_9_6# NOR2X1_34/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3875 INVX2_26/A NOR2X1_22/Y NAND2X1_26/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3876 INVX2_59/A NOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3877 vdd NOR2X1_21/Y INVX2_59/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3878 NAND2X1_25/a_9_6# NOR2X1_34/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3879 INVX2_59/A NOR2X1_21/Y NAND2X1_25/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3880 OAI21X1_60/a_9_54# INVX2_71/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3881 OAI21X1_60/Y OR2X2_0/Y OAI21X1_60/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3882 vdd OAI21X1_60/C OAI21X1_60/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3883 gnd INVX2_71/A OAI21X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3884 OAI21X1_60/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3885 OAI21X1_60/Y OAI21X1_60/C OAI21X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3886 INVX2_73/A NOR2X1_35/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3887 vdd NOR2X1_22/Y INVX2_73/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3888 NAND2X1_23/a_9_6# NOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3889 INVX2_73/A NOR2X1_22/Y NAND2X1_23/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3890 INVX2_75/A NOR2X1_35/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3891 vdd NOR2X1_21/Y INVX2_75/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3892 NAND2X1_22/a_9_6# NOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3893 INVX2_75/A NOR2X1_21/Y NAND2X1_22/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3894 INVX2_80/Y INVX2_80/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3895 INVX2_80/Y INVX2_80/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3896 vdd con_count[0] AOI22X1_60/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3897 AOI22X1_60/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3898 INVX2_80/A INVX2_126/A AOI22X1_60/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3899 AOI22X1_60/a_2_54# AOI22X1_60/C INVX2_80/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3900 AOI22X1_60/a_11_6# con_count[0] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3901 INVX2_80/A INVX2_126/Y AOI22X1_60/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3902 AOI22X1_60/a_28_6# INVX2_126/A INVX2_80/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3903 gnd AOI22X1_60/C AOI22X1_60/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3904 vdd con_count[8] AOI22X1_59/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3905 AOI22X1_59/a_2_54# INVX2_126/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3906 INVX2_79/A INVX2_126/A AOI22X1_59/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3907 AOI22X1_59/a_2_54# AOI22X1_59/C INVX2_79/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3908 AOI22X1_59/a_11_6# con_count[8] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3909 INVX2_79/A INVX2_126/Y AOI22X1_59/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3910 AOI22X1_59/a_28_6# INVX2_126/A INVX2_79/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3911 gnd AOI22X1_59/C AOI22X1_59/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3912 INVX2_79/Y INVX2_79/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3913 INVX2_79/Y INVX2_79/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3914 OAI21X1_59/a_9_54# INVX2_68/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3915 OAI21X1_59/Y OAI21X1_59/B OAI21X1_59/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3916 vdd OAI21X1_59/C OAI21X1_59/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3917 gnd INVX2_68/Y OAI21X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3918 OAI21X1_59/a_2_6# OAI21X1_59/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3919 OAI21X1_59/Y OAI21X1_59/C OAI21X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3920 vdd INVX2_43/Y DFFPOSX1_54/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3921 DFFPOSX1_54/a_17_74# OAI21X1_59/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3922 DFFPOSX1_54/a_22_6# INVX2_43/Y DFFPOSX1_54/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M3923 DFFPOSX1_54/a_31_74# DFFPOSX1_54/a_2_6# DFFPOSX1_54/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M3924 vdd DFFPOSX1_54/a_34_4# DFFPOSX1_54/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3925 DFFPOSX1_54/a_34_4# DFFPOSX1_54/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3926 DFFPOSX1_54/a_61_74# DFFPOSX1_54/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3927 DFFPOSX1_54/a_66_6# DFFPOSX1_54/a_2_6# DFFPOSX1_54/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M3928 DFFPOSX1_54/a_76_84# INVX2_43/Y DFFPOSX1_54/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3929 vdd out_win DFFPOSX1_54/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3930 gnd INVX2_43/Y DFFPOSX1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3931 out_win DFFPOSX1_54/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3932 DFFPOSX1_54/a_17_6# OAI21X1_59/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3933 DFFPOSX1_54/a_22_6# DFFPOSX1_54/a_2_6# DFFPOSX1_54/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3934 DFFPOSX1_54/a_31_6# INVX2_43/Y DFFPOSX1_54/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3935 gnd DFFPOSX1_54/a_34_4# DFFPOSX1_54/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3936 DFFPOSX1_54/a_34_4# DFFPOSX1_54/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M3937 DFFPOSX1_54/a_61_6# DFFPOSX1_54/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3938 DFFPOSX1_54/a_66_6# INVX2_43/Y DFFPOSX1_54/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M3939 DFFPOSX1_54/a_76_6# DFFPOSX1_54/a_2_6# DFFPOSX1_54/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M3940 gnd out_win DFFPOSX1_54/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3941 out_win DFFPOSX1_54/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3942 OAI21X1_58/a_9_54# AOI22X1_58/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3943 OAI21X1_58/Y XNOR2X1_41/Y OAI21X1_58/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3944 vdd NAND2X1_28/Y OAI21X1_58/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3945 gnd AOI22X1_58/Y OAI21X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3946 OAI21X1_58/a_2_6# XNOR2X1_41/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3947 OAI21X1_58/Y NAND2X1_28/Y OAI21X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3948 OAI21X1_57/a_9_54# AOI22X1_58/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3949 XOR2X1_65/A XNOR2X1_41/Y OAI21X1_57/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M3950 vdd OAI21X1_57/C XOR2X1_65/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3951 gnd AOI22X1_58/Y OAI21X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M3952 OAI21X1_57/a_2_6# XNOR2X1_41/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3953 XOR2X1_65/A OAI21X1_57/C OAI21X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3954 vdd out_MuxData[8] AOI22X1_58/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3955 AOI22X1_58/a_2_54# out_MuxData[14] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3956 AOI22X1_58/Y out_MuxData[2] AOI22X1_58/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3957 AOI22X1_58/a_2_54# XOR2X1_53/Y AOI22X1_58/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3958 AOI22X1_58/a_11_6# out_MuxData[8] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3959 AOI22X1_58/Y out_MuxData[14] AOI22X1_58/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3960 AOI22X1_58/a_28_6# out_MuxData[2] AOI22X1_58/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3961 gnd XOR2X1_53/Y AOI22X1_58/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3962 vdd INVX2_28/Y XNOR2X1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3963 XNOR2X1_36/a_18_54# XNOR2X1_36/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3964 XOR2X1_64/B XNOR2X1_36/a_2_6# XNOR2X1_36/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3965 XNOR2X1_36/a_35_54# INVX2_28/Y XOR2X1_64/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3966 vdd XOR2X1_56/Y XNOR2X1_36/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3967 XNOR2X1_36/a_12_41# XOR2X1_56/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3968 gnd INVX2_28/Y XNOR2X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3969 XNOR2X1_36/a_18_6# XNOR2X1_36/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3970 XOR2X1_64/B INVX2_28/Y XNOR2X1_36/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3971 XNOR2X1_36/a_35_6# XNOR2X1_36/a_2_6# XOR2X1_64/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3972 gnd XOR2X1_56/Y XNOR2X1_36/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3973 XNOR2X1_36/a_12_41# XOR2X1_56/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3974 vdd out_MuxData[3] AOI22X1_57/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3975 AOI22X1_57/a_2_54# out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3976 NOR2X1_28/B out_MuxData[14] AOI22X1_57/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3977 AOI22X1_57/a_2_54# XOR2X1_56/Y NOR2X1_28/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3978 AOI22X1_57/a_11_6# out_MuxData[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3979 NOR2X1_28/B out_MuxData[2] AOI22X1_57/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3980 AOI22X1_57/a_28_6# out_MuxData[14] NOR2X1_28/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3981 gnd XOR2X1_56/Y AOI22X1_57/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3982 vdd XOR2X1_57/A XOR2X1_57/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M3983 XOR2X1_57/a_18_54# XOR2X1_57/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3984 XOR2X1_57/Y XOR2X1_57/A XOR2X1_57/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M3985 XOR2X1_57/a_35_54# XOR2X1_57/a_2_6# XOR2X1_57/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M3986 vdd NOR2X1_28/Y XOR2X1_57/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3987 XOR2X1_57/a_13_43# NOR2X1_28/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M3988 gnd XOR2X1_57/A XOR2X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M3989 XOR2X1_57/a_18_6# XOR2X1_57/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3990 XOR2X1_57/Y XOR2X1_57/a_2_6# XOR2X1_57/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M3991 XOR2X1_57/a_35_6# XOR2X1_57/A XOR2X1_57/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3992 gnd NOR2X1_28/Y XOR2X1_57/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3993 XOR2X1_57/a_13_43# NOR2X1_28/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M3994 vdd XOR2X1_55/Y AOI22X1_56/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M3995 AOI22X1_56/a_2_54# INVX2_75/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3996 AND2X2_21/A INVX2_73/Y AOI22X1_56/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M3997 AOI22X1_56/a_2_54# XOR2X1_63/Y AND2X2_21/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3998 AOI22X1_56/a_11_6# XOR2X1_55/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M3999 AND2X2_21/A INVX2_75/Y AOI22X1_56/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4000 AOI22X1_56/a_28_6# INVX2_73/Y AND2X2_21/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4001 gnd XOR2X1_63/Y AOI22X1_56/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4002 vdd XOR2X1_55/A XOR2X1_55/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4003 XOR2X1_55/a_18_54# XOR2X1_55/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4004 XOR2X1_55/Y XOR2X1_55/A XOR2X1_55/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4005 XOR2X1_55/a_35_54# XOR2X1_55/a_2_6# XOR2X1_55/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4006 vdd XOR2X1_55/B XOR2X1_55/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4007 XOR2X1_55/a_13_43# XOR2X1_55/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4008 gnd XOR2X1_55/A XOR2X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4009 XOR2X1_55/a_18_6# XOR2X1_55/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4010 XOR2X1_55/Y XOR2X1_55/a_2_6# XOR2X1_55/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4011 XOR2X1_55/a_35_6# XOR2X1_55/A XOR2X1_55/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4012 gnd XOR2X1_55/B XOR2X1_55/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4013 XOR2X1_55/a_13_43# XOR2X1_55/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4014 NAND3X1_25/Y XOR2X1_55/B vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4015 vdd NAND3X1_25/B NAND3X1_25/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4016 NAND3X1_25/Y XOR2X1_55/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4017 NAND3X1_25/a_9_6# XOR2X1_55/B gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4018 NAND3X1_25/a_14_6# NAND3X1_25/B NAND3X1_25/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4019 NAND3X1_25/Y XOR2X1_55/A NAND3X1_25/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4020 vdd NOR2X1_27/A AOI21X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M4021 AOI21X1_6/a_2_54# AOI21X1_6/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4022 INVX2_67/A NOR2X1_27/Y AOI21X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4023 AOI21X1_6/a_12_6# NOR2X1_27/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4024 INVX2_67/A AOI21X1_6/B AOI21X1_6/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M4025 gnd NOR2X1_27/Y INVX2_67/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4026 vdd out_MuxData[2] AOI22X1_54/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4027 AOI22X1_54/a_2_54# out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4028 NOR2X1_27/A out_MuxData[13] AOI22X1_54/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4029 AOI22X1_54/a_2_54# XOR2X1_60/Y NOR2X1_27/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4030 AOI22X1_54/a_11_6# out_MuxData[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4031 NOR2X1_27/A out_MuxData[1] AOI22X1_54/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4032 AOI22X1_54/a_28_6# out_MuxData[13] NOR2X1_27/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4033 gnd XOR2X1_60/Y AOI22X1_54/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4034 OAI22X1_9/a_9_54# INVX2_65/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4035 OAI22X1_9/Y INVX2_84/Y OAI22X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4036 OAI22X1_9/a_28_54# INVX2_99/Y OAI22X1_9/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4037 vdd INVX2_85/Y OAI22X1_9/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4038 gnd INVX2_65/Y OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4039 OAI22X1_9/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4040 OAI22X1_9/Y INVX2_99/Y OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4041 OAI22X1_9/a_2_6# INVX2_85/Y OAI22X1_9/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4042 vdd BUFX2_5/Y DFFPOSX1_52/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4043 DFFPOSX1_52/a_17_74# INVX2_78/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4044 DFFPOSX1_52/a_22_6# BUFX2_5/Y DFFPOSX1_52/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4045 DFFPOSX1_52/a_31_74# DFFPOSX1_52/a_2_6# DFFPOSX1_52/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4046 vdd DFFPOSX1_52/a_34_4# DFFPOSX1_52/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4047 DFFPOSX1_52/a_34_4# DFFPOSX1_52/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4048 DFFPOSX1_52/a_61_74# DFFPOSX1_52/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4049 DFFPOSX1_52/a_66_6# DFFPOSX1_52/a_2_6# DFFPOSX1_52/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4050 DFFPOSX1_52/a_76_84# BUFX2_5/Y DFFPOSX1_52/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4051 vdd out_MuxData[14] DFFPOSX1_52/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4052 gnd BUFX2_5/Y DFFPOSX1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4053 out_MuxData[14] DFFPOSX1_52/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4054 DFFPOSX1_52/a_17_6# INVX2_78/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4055 DFFPOSX1_52/a_22_6# DFFPOSX1_52/a_2_6# DFFPOSX1_52/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4056 DFFPOSX1_52/a_31_6# BUFX2_5/Y DFFPOSX1_52/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4057 gnd DFFPOSX1_52/a_34_4# DFFPOSX1_52/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4058 DFFPOSX1_52/a_34_4# DFFPOSX1_52/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4059 DFFPOSX1_52/a_61_6# DFFPOSX1_52/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4060 DFFPOSX1_52/a_66_6# BUFX2_5/Y DFFPOSX1_52/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4061 DFFPOSX1_52/a_76_6# DFFPOSX1_52/a_2_6# DFFPOSX1_52/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4062 gnd out_MuxData[14] DFFPOSX1_52/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4063 out_MuxData[14] DFFPOSX1_52/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4064 INVX2_78/Y INVX2_78/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4065 INVX2_78/Y INVX2_78/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4066 vdd AOI22X1_51/B AOI22X1_53/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4067 AOI22X1_53/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4068 INVX2_78/A INVX2_99/A AOI22X1_53/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4069 AOI22X1_53/a_2_54# out_MuxData[14] INVX2_78/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4070 AOI22X1_53/a_11_6# AOI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4071 INVX2_78/A con_writeout AOI22X1_53/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4072 AOI22X1_53/a_28_6# INVX2_99/A INVX2_78/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4073 gnd out_MuxData[14] AOI22X1_53/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4074 vdd INVX2_61/Y DFFPOSX1_50/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4075 DFFPOSX1_50/a_17_74# INVX2_76/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4076 DFFPOSX1_50/a_22_6# INVX2_61/Y DFFPOSX1_50/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4077 DFFPOSX1_50/a_31_74# DFFPOSX1_50/a_2_6# DFFPOSX1_50/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4078 vdd DFFPOSX1_50/a_34_4# DFFPOSX1_50/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4079 DFFPOSX1_50/a_34_4# DFFPOSX1_50/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4080 DFFPOSX1_50/a_61_74# DFFPOSX1_50/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4081 DFFPOSX1_50/a_66_6# DFFPOSX1_50/a_2_6# DFFPOSX1_50/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4082 DFFPOSX1_50/a_76_84# INVX2_61/Y DFFPOSX1_50/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4083 vdd AOI22X1_51/B DFFPOSX1_50/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4084 gnd INVX2_61/Y DFFPOSX1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4085 AOI22X1_51/B DFFPOSX1_50/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4086 DFFPOSX1_50/a_17_6# INVX2_76/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4087 DFFPOSX1_50/a_22_6# DFFPOSX1_50/a_2_6# DFFPOSX1_50/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4088 DFFPOSX1_50/a_31_6# INVX2_61/Y DFFPOSX1_50/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4089 gnd DFFPOSX1_50/a_34_4# DFFPOSX1_50/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4090 DFFPOSX1_50/a_34_4# DFFPOSX1_50/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4091 DFFPOSX1_50/a_61_6# DFFPOSX1_50/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4092 DFFPOSX1_50/a_66_6# INVX2_61/Y DFFPOSX1_50/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4093 DFFPOSX1_50/a_76_6# DFFPOSX1_50/a_2_6# DFFPOSX1_50/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4094 gnd AOI22X1_51/B DFFPOSX1_50/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4095 AOI22X1_51/B DFFPOSX1_50/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4096 INVX2_77/Y INVX2_77/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4097 INVX2_77/Y INVX2_77/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4098 INVX2_76/Y INVX2_76/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4099 INVX2_76/Y INVX2_76/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4100 vdd con_restart AOI22X1_51/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4101 AOI22X1_51/a_2_54# AOI22X1_51/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4102 INVX2_76/A out_MemBData[14] AOI22X1_51/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4103 AOI22X1_51/a_2_54# BUFX2_7/Y INVX2_76/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4104 AOI22X1_51/a_11_6# con_restart gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4105 INVX2_76/A AOI22X1_51/B AOI22X1_51/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4106 AOI22X1_51/a_28_6# out_MemBData[14] INVX2_76/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4107 gnd BUFX2_7/Y AOI22X1_51/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4108 vdd BUFX2_8/A BUFX2_8/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4109 BUFX2_8/Y BUFX2_8/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4110 gnd BUFX2_8/A BUFX2_8/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4111 BUFX2_8/Y BUFX2_8/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4112 INVX2_75/Y INVX2_75/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4113 INVX2_75/Y INVX2_75/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4114 INVX2_73/Y INVX2_73/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4115 INVX2_73/Y INVX2_73/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4116 vdd BUFX2_5/Y DFFPOSX1_48/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4117 DFFPOSX1_48/a_17_74# OAI21X1_61/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4118 DFFPOSX1_48/a_22_6# BUFX2_5/Y DFFPOSX1_48/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4119 DFFPOSX1_48/a_31_74# DFFPOSX1_48/a_2_6# DFFPOSX1_48/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4120 vdd DFFPOSX1_48/a_34_4# DFFPOSX1_48/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4121 DFFPOSX1_48/a_34_4# DFFPOSX1_48/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4122 DFFPOSX1_48/a_61_74# DFFPOSX1_48/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4123 DFFPOSX1_48/a_66_6# DFFPOSX1_48/a_2_6# DFFPOSX1_48/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4124 DFFPOSX1_48/a_76_84# BUFX2_5/Y DFFPOSX1_48/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4125 vdd out_MemBData[14] DFFPOSX1_48/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4126 gnd BUFX2_5/Y DFFPOSX1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4127 out_MemBData[14] DFFPOSX1_48/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4128 DFFPOSX1_48/a_17_6# OAI21X1_61/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4129 DFFPOSX1_48/a_22_6# DFFPOSX1_48/a_2_6# DFFPOSX1_48/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4130 DFFPOSX1_48/a_31_6# BUFX2_5/Y DFFPOSX1_48/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4131 gnd DFFPOSX1_48/a_34_4# DFFPOSX1_48/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4132 DFFPOSX1_48/a_34_4# DFFPOSX1_48/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4133 DFFPOSX1_48/a_61_6# DFFPOSX1_48/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4134 DFFPOSX1_48/a_66_6# BUFX2_5/Y DFFPOSX1_48/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4135 DFFPOSX1_48/a_76_6# DFFPOSX1_48/a_2_6# DFFPOSX1_48/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4136 gnd out_MemBData[14] DFFPOSX1_48/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4137 out_MemBData[14] DFFPOSX1_48/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4138 OAI21X1_53/a_9_54# NOR2X1_19/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4139 OAI21X1_60/C AND2X2_19/Y OAI21X1_53/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4140 vdd out_MemBData[0] OAI21X1_60/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4141 gnd NOR2X1_19/Y OAI21X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4142 OAI21X1_53/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4143 OAI21X1_60/C out_MemBData[0] OAI21X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4144 vdd BUFX2_6/Y DFFPOSX1_46/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4145 DFFPOSX1_46/a_17_74# OAI21X1_60/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4146 DFFPOSX1_46/a_22_6# BUFX2_6/Y DFFPOSX1_46/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4147 DFFPOSX1_46/a_31_74# DFFPOSX1_46/a_2_6# DFFPOSX1_46/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4148 vdd DFFPOSX1_46/a_34_4# DFFPOSX1_46/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4149 DFFPOSX1_46/a_34_4# DFFPOSX1_46/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4150 DFFPOSX1_46/a_61_74# DFFPOSX1_46/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4151 DFFPOSX1_46/a_66_6# DFFPOSX1_46/a_2_6# DFFPOSX1_46/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4152 DFFPOSX1_46/a_76_84# BUFX2_6/Y DFFPOSX1_46/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4153 vdd out_MemBData[0] DFFPOSX1_46/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4154 gnd BUFX2_6/Y DFFPOSX1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4155 out_MemBData[0] DFFPOSX1_46/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4156 DFFPOSX1_46/a_17_6# OAI21X1_60/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4157 DFFPOSX1_46/a_22_6# DFFPOSX1_46/a_2_6# DFFPOSX1_46/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4158 DFFPOSX1_46/a_31_6# BUFX2_6/Y DFFPOSX1_46/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4159 gnd DFFPOSX1_46/a_34_4# DFFPOSX1_46/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4160 DFFPOSX1_46/a_34_4# DFFPOSX1_46/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4161 DFFPOSX1_46/a_61_6# DFFPOSX1_46/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4162 DFFPOSX1_46/a_66_6# BUFX2_6/Y DFFPOSX1_46/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4163 DFFPOSX1_46/a_76_6# DFFPOSX1_46/a_2_6# DFFPOSX1_46/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4164 gnd out_MemBData[0] DFFPOSX1_46/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4165 out_MemBData[0] DFFPOSX1_46/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4166 vdd in_clka BUFX2_6/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4167 BUFX2_6/Y BUFX2_6/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4168 gnd in_clka BUFX2_6/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4169 BUFX2_6/Y BUFX2_6/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4170 vdd in_clka BUFX2_5/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4171 BUFX2_5/Y BUFX2_5/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4172 gnd in_clka BUFX2_5/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4173 BUFX2_5/Y BUFX2_5/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4174 vdd INVX2_41/Y DFFPOSX1_45/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4175 DFFPOSX1_45/a_17_74# INVX2_80/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4176 DFFPOSX1_45/a_22_6# INVX2_41/Y DFFPOSX1_45/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4177 DFFPOSX1_45/a_31_74# DFFPOSX1_45/a_2_6# DFFPOSX1_45/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4178 vdd DFFPOSX1_45/a_34_4# DFFPOSX1_45/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4179 DFFPOSX1_45/a_34_4# DFFPOSX1_45/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4180 DFFPOSX1_45/a_61_74# DFFPOSX1_45/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4181 DFFPOSX1_45/a_66_6# DFFPOSX1_45/a_2_6# DFFPOSX1_45/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4182 DFFPOSX1_45/a_76_84# INVX2_41/Y DFFPOSX1_45/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4183 vdd con_count[0] DFFPOSX1_45/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4184 gnd INVX2_41/Y DFFPOSX1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4185 con_count[0] DFFPOSX1_45/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4186 DFFPOSX1_45/a_17_6# INVX2_80/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4187 DFFPOSX1_45/a_22_6# DFFPOSX1_45/a_2_6# DFFPOSX1_45/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4188 DFFPOSX1_45/a_31_6# INVX2_41/Y DFFPOSX1_45/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4189 gnd DFFPOSX1_45/a_34_4# DFFPOSX1_45/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4190 DFFPOSX1_45/a_34_4# DFFPOSX1_45/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4191 DFFPOSX1_45/a_61_6# DFFPOSX1_45/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4192 DFFPOSX1_45/a_66_6# INVX2_41/Y DFFPOSX1_45/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4193 DFFPOSX1_45/a_76_6# DFFPOSX1_45/a_2_6# DFFPOSX1_45/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4194 gnd con_count[0] DFFPOSX1_45/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4195 con_count[0] DFFPOSX1_45/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4196 INVX2_72/Y INVX2_72/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4197 INVX2_72/Y INVX2_72/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4198 INVX2_126/A OAI21X1_52/C vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4199 vdd INVX2_53/A INVX2_126/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4200 NAND2X1_21/a_9_6# OAI21X1_52/C gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4201 INVX2_126/A INVX2_53/A NAND2X1_21/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4202 vdd INVX2_41/Y DFFPOSX1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4203 DFFPOSX1_42/a_17_74# INVX2_79/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4204 DFFPOSX1_42/a_22_6# INVX2_41/Y DFFPOSX1_42/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4205 DFFPOSX1_42/a_31_74# DFFPOSX1_42/a_2_6# DFFPOSX1_42/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4206 vdd DFFPOSX1_42/a_34_4# DFFPOSX1_42/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4207 DFFPOSX1_42/a_34_4# DFFPOSX1_42/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4208 DFFPOSX1_42/a_61_74# DFFPOSX1_42/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4209 DFFPOSX1_42/a_66_6# DFFPOSX1_42/a_2_6# DFFPOSX1_42/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4210 DFFPOSX1_42/a_76_84# INVX2_41/Y DFFPOSX1_42/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4211 vdd con_count[8] DFFPOSX1_42/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4212 gnd INVX2_41/Y DFFPOSX1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4213 con_count[8] DFFPOSX1_42/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4214 DFFPOSX1_42/a_17_6# INVX2_79/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4215 DFFPOSX1_42/a_22_6# DFFPOSX1_42/a_2_6# DFFPOSX1_42/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4216 DFFPOSX1_42/a_31_6# INVX2_41/Y DFFPOSX1_42/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4217 gnd DFFPOSX1_42/a_34_4# DFFPOSX1_42/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4218 DFFPOSX1_42/a_34_4# DFFPOSX1_42/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4219 DFFPOSX1_42/a_61_6# DFFPOSX1_42/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4220 DFFPOSX1_42/a_66_6# INVX2_41/Y DFFPOSX1_42/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4221 DFFPOSX1_42/a_76_6# DFFPOSX1_42/a_2_6# DFFPOSX1_42/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4222 gnd con_count[8] DFFPOSX1_42/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4223 con_count[8] DFFPOSX1_42/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4224 OAI21X1_52/a_9_54# INVX2_51/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4225 OAI21X1_59/B INVX2_52/Y OAI21X1_52/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4226 vdd OAI21X1_52/C OAI21X1_59/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4227 gnd INVX2_51/A OAI21X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4228 OAI21X1_52/a_2_6# INVX2_52/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4229 OAI21X1_59/B OAI21X1_52/C OAI21X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4230 INVX2_68/Y out_win vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4231 INVX2_68/Y out_win gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4232 AND2X2_24/a_2_6# XOR2X1_58/B vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4233 vdd XOR2X1_58/A AND2X2_24/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4234 AND2X2_24/Y AND2X2_24/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4235 AND2X2_24/a_9_6# XOR2X1_58/B AND2X2_24/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4236 gnd XOR2X1_58/A AND2X2_24/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4237 AND2X2_24/Y AND2X2_24/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4238 OAI21X1_57/C XOR2X1_58/B vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4239 vdd NAND2X1_28/Y OAI21X1_57/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4240 OAI21X1_57/C XOR2X1_58/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4241 NAND3X1_26/a_9_6# XOR2X1_58/B gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4242 NAND3X1_26/a_14_6# NAND2X1_28/Y NAND3X1_26/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4243 OAI21X1_57/C XOR2X1_58/A NAND3X1_26/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4244 vdd XOR2X1_58/A XOR2X1_58/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4245 XOR2X1_58/a_18_54# XOR2X1_58/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4246 XOR2X1_58/Y XOR2X1_58/A XOR2X1_58/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4247 XOR2X1_58/a_35_54# XOR2X1_58/a_2_6# XOR2X1_58/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4248 vdd XOR2X1_58/B XOR2X1_58/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4249 XOR2X1_58/a_13_43# XOR2X1_58/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4250 gnd XOR2X1_58/A XOR2X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4251 XOR2X1_58/a_18_6# XOR2X1_58/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4252 XOR2X1_58/Y XOR2X1_58/a_2_6# XOR2X1_58/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4253 XOR2X1_58/a_35_6# XOR2X1_58/A XOR2X1_58/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4254 gnd XOR2X1_58/B XOR2X1_58/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4255 XOR2X1_58/a_13_43# XOR2X1_58/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4256 vdd INVX2_85/Y XNOR2X1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4257 XNOR2X1_35/a_18_54# XNOR2X1_35/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4258 XOR2X1_58/A XNOR2X1_35/a_2_6# XNOR2X1_35/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4259 XNOR2X1_35/a_35_54# INVX2_85/Y XOR2X1_58/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4260 vdd XOR2X1_53/Y XNOR2X1_35/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4261 XNOR2X1_35/a_12_41# XOR2X1_53/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4262 gnd INVX2_85/Y XNOR2X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4263 XNOR2X1_35/a_18_6# XNOR2X1_35/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4264 XOR2X1_58/A INVX2_85/Y XNOR2X1_35/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4265 XNOR2X1_35/a_35_6# XNOR2X1_35/a_2_6# XOR2X1_58/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4266 gnd XOR2X1_53/Y XNOR2X1_35/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4267 XNOR2X1_35/a_12_41# XOR2X1_53/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4268 vdd INVX2_85/Y XOR2X1_56/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4269 XOR2X1_56/a_18_54# XOR2X1_56/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4270 XOR2X1_56/Y INVX2_85/Y XOR2X1_56/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4271 XOR2X1_56/a_35_54# XOR2X1_56/a_2_6# XOR2X1_56/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4272 vdd INVX2_86/Y XOR2X1_56/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4273 XOR2X1_56/a_13_43# INVX2_86/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4274 gnd INVX2_85/Y XOR2X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4275 XOR2X1_56/a_18_6# XOR2X1_56/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4276 XOR2X1_56/Y XOR2X1_56/a_2_6# XOR2X1_56/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4277 XOR2X1_56/a_35_6# INVX2_85/Y XOR2X1_56/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4278 gnd INVX2_86/Y XOR2X1_56/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4279 XOR2X1_56/a_13_43# INVX2_86/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4280 vdd INVX2_73/Y AOI22X1_55/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4281 AOI22X1_55/a_2_54# XNOR2X1_45/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4282 AOI22X1_55/Y AOI22X1_55/D AOI22X1_55/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4283 AOI22X1_55/a_2_54# INVX2_75/Y AOI22X1_55/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4284 AOI22X1_55/a_11_6# INVX2_73/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4285 AOI22X1_55/Y XNOR2X1_45/Y AOI22X1_55/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4286 AOI22X1_55/a_28_6# AOI22X1_55/D AOI22X1_55/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4287 gnd INVX2_75/Y AOI22X1_55/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4288 AND2X2_23/a_2_6# XOR2X1_55/B vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4289 vdd XOR2X1_55/A AND2X2_23/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4290 AND2X2_23/Y AND2X2_23/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4291 AND2X2_23/a_9_6# XOR2X1_55/B AND2X2_23/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4292 gnd XOR2X1_55/A AND2X2_23/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4293 AND2X2_23/Y AND2X2_23/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4294 OAI21X1_56/a_9_54# OAI21X1_56/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4295 XOR2X1_61/A INVX2_67/Y OAI21X1_56/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4296 vdd NAND3X1_25/Y XOR2X1_61/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4297 gnd OAI21X1_56/A OAI21X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4298 OAI21X1_56/a_2_6# INVX2_67/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4299 XOR2X1_61/A NAND3X1_25/Y OAI21X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4300 vdd BUFX2_11/Y DFFPOSX1_53/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4301 DFFPOSX1_53/a_17_74# OAI22X1_9/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4302 DFFPOSX1_53/a_22_6# BUFX2_11/Y DFFPOSX1_53/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4303 DFFPOSX1_53/a_31_74# DFFPOSX1_53/a_2_6# DFFPOSX1_53/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4304 vdd DFFPOSX1_53/a_34_4# DFFPOSX1_53/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4305 DFFPOSX1_53/a_34_4# DFFPOSX1_53/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4306 DFFPOSX1_53/a_61_74# DFFPOSX1_53/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4307 DFFPOSX1_53/a_66_6# DFFPOSX1_53/a_2_6# DFFPOSX1_53/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4308 DFFPOSX1_53/a_76_84# BUFX2_11/Y DFFPOSX1_53/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4309 vdd out_MuxData[2] DFFPOSX1_53/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4310 gnd BUFX2_11/Y DFFPOSX1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4311 out_MuxData[2] DFFPOSX1_53/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4312 DFFPOSX1_53/a_17_6# OAI22X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4313 DFFPOSX1_53/a_22_6# DFFPOSX1_53/a_2_6# DFFPOSX1_53/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4314 DFFPOSX1_53/a_31_6# BUFX2_11/Y DFFPOSX1_53/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4315 gnd DFFPOSX1_53/a_34_4# DFFPOSX1_53/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4316 DFFPOSX1_53/a_34_4# DFFPOSX1_53/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4317 DFFPOSX1_53/a_61_6# DFFPOSX1_53/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4318 DFFPOSX1_53/a_66_6# BUFX2_11/Y DFFPOSX1_53/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4319 DFFPOSX1_53/a_76_6# DFFPOSX1_53/a_2_6# DFFPOSX1_53/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4320 gnd out_MuxData[2] DFFPOSX1_53/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4321 out_MuxData[2] DFFPOSX1_53/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4322 vdd BUFX2_5/Y DFFPOSX1_51/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4323 DFFPOSX1_51/a_17_74# OAI22X1_6/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4324 DFFPOSX1_51/a_22_6# BUFX2_5/Y DFFPOSX1_51/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4325 DFFPOSX1_51/a_31_74# DFFPOSX1_51/a_2_6# DFFPOSX1_51/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4326 vdd DFFPOSX1_51/a_34_4# DFFPOSX1_51/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4327 DFFPOSX1_51/a_34_4# DFFPOSX1_51/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4328 DFFPOSX1_51/a_61_74# DFFPOSX1_51/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4329 DFFPOSX1_51/a_66_6# DFFPOSX1_51/a_2_6# DFFPOSX1_51/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4330 DFFPOSX1_51/a_76_84# BUFX2_5/Y DFFPOSX1_51/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4331 vdd out_MuxData[0] DFFPOSX1_51/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4332 gnd BUFX2_5/Y DFFPOSX1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4333 out_MuxData[0] DFFPOSX1_51/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4334 DFFPOSX1_51/a_17_6# OAI22X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4335 DFFPOSX1_51/a_22_6# DFFPOSX1_51/a_2_6# DFFPOSX1_51/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4336 DFFPOSX1_51/a_31_6# BUFX2_5/Y DFFPOSX1_51/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4337 gnd DFFPOSX1_51/a_34_4# DFFPOSX1_51/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4338 DFFPOSX1_51/a_34_4# DFFPOSX1_51/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4339 DFFPOSX1_51/a_61_6# DFFPOSX1_51/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4340 DFFPOSX1_51/a_66_6# BUFX2_5/Y DFFPOSX1_51/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4341 DFFPOSX1_51/a_76_6# DFFPOSX1_51/a_2_6# DFFPOSX1_51/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4342 gnd out_MuxData[0] DFFPOSX1_51/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4343 out_MuxData[0] DFFPOSX1_51/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4344 vdd AOI22X1_50/B AOI22X1_52/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4345 AOI22X1_52/a_2_54# con_writeout vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4346 INVX2_66/A INVX2_99/A AOI22X1_52/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4347 AOI22X1_52/a_2_54# out_MuxData[15] INVX2_66/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4348 AOI22X1_52/a_11_6# AOI22X1_50/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4349 INVX2_66/A con_writeout AOI22X1_52/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4350 AOI22X1_52/a_28_6# INVX2_99/A INVX2_66/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4351 gnd out_MuxData[15] AOI22X1_52/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4352 vdd INVX2_61/Y DFFPOSX1_49/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4353 DFFPOSX1_49/a_17_74# INVX2_77/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4354 DFFPOSX1_49/a_22_6# INVX2_61/Y DFFPOSX1_49/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4355 DFFPOSX1_49/a_31_74# DFFPOSX1_49/a_2_6# DFFPOSX1_49/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4356 vdd DFFPOSX1_49/a_34_4# DFFPOSX1_49/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4357 DFFPOSX1_49/a_34_4# DFFPOSX1_49/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4358 DFFPOSX1_49/a_61_74# DFFPOSX1_49/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4359 DFFPOSX1_49/a_66_6# DFFPOSX1_49/a_2_6# DFFPOSX1_49/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4360 DFFPOSX1_49/a_76_84# INVX2_61/Y DFFPOSX1_49/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4361 vdd AOI22X1_50/B DFFPOSX1_49/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4362 gnd INVX2_61/Y DFFPOSX1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4363 AOI22X1_50/B DFFPOSX1_49/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4364 DFFPOSX1_49/a_17_6# INVX2_77/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4365 DFFPOSX1_49/a_22_6# DFFPOSX1_49/a_2_6# DFFPOSX1_49/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4366 DFFPOSX1_49/a_31_6# INVX2_61/Y DFFPOSX1_49/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4367 gnd DFFPOSX1_49/a_34_4# DFFPOSX1_49/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4368 DFFPOSX1_49/a_34_4# DFFPOSX1_49/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4369 DFFPOSX1_49/a_61_6# DFFPOSX1_49/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4370 DFFPOSX1_49/a_66_6# INVX2_61/Y DFFPOSX1_49/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4371 DFFPOSX1_49/a_76_6# DFFPOSX1_49/a_2_6# DFFPOSX1_49/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4372 gnd AOI22X1_50/B DFFPOSX1_49/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4373 AOI22X1_50/B DFFPOSX1_49/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4374 vdd con_restart AOI22X1_50/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4375 AOI22X1_50/a_2_54# AOI22X1_50/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4376 INVX2_77/A out_MemBData[15] AOI22X1_50/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4377 AOI22X1_50/a_2_54# BUFX2_7/Y INVX2_77/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4378 AOI22X1_50/a_11_6# con_restart gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4379 INVX2_77/A AOI22X1_50/B AOI22X1_50/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4380 AOI22X1_50/a_28_6# out_MemBData[15] INVX2_77/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4381 gnd BUFX2_7/Y AOI22X1_50/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4382 vdd BUFX2_8/A BUFX2_7/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4383 BUFX2_7/Y BUFX2_7/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4384 gnd BUFX2_8/A BUFX2_7/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4385 BUFX2_7/Y BUFX2_7/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4386 BUFX2_8/A con_restart vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4387 BUFX2_8/A con_restart gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4388 NOR2X1_20/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4389 NOR2X1_20/Y INVX2_73/Y NOR2X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4390 NOR2X1_20/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M4391 gnd INVX2_73/Y NOR2X1_20/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4392 OAI21X1_55/a_9_54# NOR2X1_20/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4393 OAI21X1_55/Y AND2X2_19/Y OAI21X1_55/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4394 vdd out_MemBData[15] OAI21X1_55/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4395 gnd NOR2X1_20/Y OAI21X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4396 OAI21X1_55/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4397 OAI21X1_55/Y out_MemBData[15] OAI21X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4398 OAI21X1_54/a_9_54# INVX2_73/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4399 OAI21X1_54/Y OR2X2_0/Y OAI21X1_54/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4400 vdd OAI21X1_55/Y OAI21X1_54/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4401 gnd INVX2_73/A OAI21X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4402 OAI21X1_54/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4403 OAI21X1_54/Y OAI21X1_55/Y OAI21X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4404 vdd BUFX2_5/Y DFFPOSX1_47/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4405 DFFPOSX1_47/a_17_74# OAI21X1_54/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4406 DFFPOSX1_47/a_22_6# BUFX2_5/Y DFFPOSX1_47/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4407 DFFPOSX1_47/a_31_74# DFFPOSX1_47/a_2_6# DFFPOSX1_47/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4408 vdd DFFPOSX1_47/a_34_4# DFFPOSX1_47/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4409 DFFPOSX1_47/a_34_4# DFFPOSX1_47/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4410 DFFPOSX1_47/a_61_74# DFFPOSX1_47/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4411 DFFPOSX1_47/a_66_6# DFFPOSX1_47/a_2_6# DFFPOSX1_47/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4412 DFFPOSX1_47/a_76_84# BUFX2_5/Y DFFPOSX1_47/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4413 vdd out_MemBData[15] DFFPOSX1_47/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4414 gnd BUFX2_5/Y DFFPOSX1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4415 out_MemBData[15] DFFPOSX1_47/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4416 DFFPOSX1_47/a_17_6# OAI21X1_54/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4417 DFFPOSX1_47/a_22_6# DFFPOSX1_47/a_2_6# DFFPOSX1_47/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4418 DFFPOSX1_47/a_31_6# BUFX2_5/Y DFFPOSX1_47/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4419 gnd DFFPOSX1_47/a_34_4# DFFPOSX1_47/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4420 DFFPOSX1_47/a_34_4# DFFPOSX1_47/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4421 DFFPOSX1_47/a_61_6# DFFPOSX1_47/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4422 DFFPOSX1_47/a_66_6# BUFX2_5/Y DFFPOSX1_47/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4423 DFFPOSX1_47/a_76_6# DFFPOSX1_47/a_2_6# DFFPOSX1_47/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4424 gnd out_MemBData[15] DFFPOSX1_47/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4425 out_MemBData[15] DFFPOSX1_47/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4426 NOR2X1_19/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4427 NOR2X1_19/Y INVX2_71/Y NOR2X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4428 NOR2X1_19/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M4429 gnd INVX2_71/Y NOR2X1_19/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4430 INVX2_71/Y INVX2_71/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4431 INVX2_71/Y INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4432 vdd BUFX2_6/Y DFFPOSX1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4433 DFFPOSX1_44/a_17_74# OAI21X1_45/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4434 DFFPOSX1_44/a_22_6# BUFX2_6/Y DFFPOSX1_44/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4435 DFFPOSX1_44/a_31_74# DFFPOSX1_44/a_2_6# DFFPOSX1_44/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4436 vdd DFFPOSX1_44/a_34_4# DFFPOSX1_44/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4437 DFFPOSX1_44/a_34_4# DFFPOSX1_44/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4438 DFFPOSX1_44/a_61_74# DFFPOSX1_44/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4439 DFFPOSX1_44/a_66_6# DFFPOSX1_44/a_2_6# DFFPOSX1_44/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4440 DFFPOSX1_44/a_76_84# BUFX2_6/Y DFFPOSX1_44/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4441 vdd INVX2_57/A DFFPOSX1_44/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4442 gnd BUFX2_6/Y DFFPOSX1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4443 INVX2_57/A DFFPOSX1_44/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4444 DFFPOSX1_44/a_17_6# OAI21X1_45/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4445 DFFPOSX1_44/a_22_6# DFFPOSX1_44/a_2_6# DFFPOSX1_44/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4446 DFFPOSX1_44/a_31_6# BUFX2_6/Y DFFPOSX1_44/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4447 gnd DFFPOSX1_44/a_34_4# DFFPOSX1_44/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4448 DFFPOSX1_44/a_34_4# DFFPOSX1_44/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4449 DFFPOSX1_44/a_61_6# DFFPOSX1_44/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4450 DFFPOSX1_44/a_66_6# BUFX2_6/Y DFFPOSX1_44/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4451 DFFPOSX1_44/a_76_6# DFFPOSX1_44/a_2_6# DFFPOSX1_44/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4452 gnd INVX2_57/A DFFPOSX1_44/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4453 INVX2_57/A DFFPOSX1_44/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4454 vdd INVX2_41/Y DFFPOSX1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4455 DFFPOSX1_43/a_17_74# INVX2_69/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4456 DFFPOSX1_43/a_22_6# INVX2_41/Y DFFPOSX1_43/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4457 DFFPOSX1_43/a_31_74# DFFPOSX1_43/a_2_6# DFFPOSX1_43/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4458 vdd DFFPOSX1_43/a_34_4# DFFPOSX1_43/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4459 DFFPOSX1_43/a_34_4# DFFPOSX1_43/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4460 DFFPOSX1_43/a_61_74# DFFPOSX1_43/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4461 DFFPOSX1_43/a_66_6# DFFPOSX1_43/a_2_6# DFFPOSX1_43/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4462 DFFPOSX1_43/a_76_84# INVX2_41/Y DFFPOSX1_43/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4463 vdd con_readData DFFPOSX1_43/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4464 gnd INVX2_41/Y DFFPOSX1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4465 con_readData DFFPOSX1_43/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4466 DFFPOSX1_43/a_17_6# INVX2_69/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4467 DFFPOSX1_43/a_22_6# DFFPOSX1_43/a_2_6# DFFPOSX1_43/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4468 DFFPOSX1_43/a_31_6# INVX2_41/Y DFFPOSX1_43/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4469 gnd DFFPOSX1_43/a_34_4# DFFPOSX1_43/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4470 DFFPOSX1_43/a_34_4# DFFPOSX1_43/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4471 DFFPOSX1_43/a_61_6# DFFPOSX1_43/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4472 DFFPOSX1_43/a_66_6# INVX2_41/Y DFFPOSX1_43/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4473 DFFPOSX1_43/a_76_6# DFFPOSX1_43/a_2_6# DFFPOSX1_43/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4474 gnd con_readData DFFPOSX1_43/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4475 con_readData DFFPOSX1_43/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4476 NOR2X1_18/a_9_54# INVX2_55/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4477 INVX2_53/A INVX2_69/Y NOR2X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4478 INVX2_53/A INVX2_55/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M4479 gnd INVX2_69/Y INVX2_53/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4480 INVX2_70/Y INVX2_70/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4481 INVX2_70/Y INVX2_70/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4482 INVX2_69/Y INVX2_69/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4483 INVX2_69/Y INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4484 OAI21X1_59/C INVX2_52/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4485 vdd INVX2_40/Y OAI21X1_59/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4486 OAI21X1_59/C INVX2_51/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4487 NAND3X1_24/a_9_6# INVX2_52/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4488 NAND3X1_24/a_14_6# INVX2_40/Y NAND3X1_24/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4489 OAI21X1_59/C INVX2_51/A NAND3X1_24/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4490 INVX2_69/A INVX2_51/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4491 vdd INVX2_40/Y INVX2_69/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4492 INVX2_69/A INVX2_52/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4493 NAND3X1_23/a_9_6# INVX2_51/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4494 NAND3X1_23/a_14_6# INVX2_40/Y NAND3X1_23/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4495 INVX2_69/A INVX2_52/A NAND3X1_23/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4496 vdd OAI21X1_58/Y XNOR2X1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4497 XNOR2X1_34/a_18_54# XNOR2X1_34/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4498 AOI22X1_48/B XNOR2X1_34/a_2_6# XNOR2X1_34/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4499 XNOR2X1_34/a_35_54# OAI21X1_58/Y AOI22X1_48/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4500 vdd AND2X2_24/Y XNOR2X1_34/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4501 XNOR2X1_34/a_12_41# AND2X2_24/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4502 gnd OAI21X1_58/Y XNOR2X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4503 XNOR2X1_34/a_18_6# XNOR2X1_34/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4504 AOI22X1_48/B OAI21X1_58/Y XNOR2X1_34/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4505 XNOR2X1_34/a_35_6# XNOR2X1_34/a_2_6# AOI22X1_48/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4506 gnd AND2X2_24/Y XNOR2X1_34/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4507 XNOR2X1_34/a_12_41# AND2X2_24/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4508 vdd OAI21X1_51/Y XNOR2X1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4509 XNOR2X1_33/a_18_54# XNOR2X1_33/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4510 AOI22X1_48/D XNOR2X1_33/a_2_6# XNOR2X1_33/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4511 XNOR2X1_33/a_35_54# OAI21X1_51/Y AOI22X1_48/D vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4512 vdd AND2X2_22/Y XNOR2X1_33/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4513 XNOR2X1_33/a_12_41# AND2X2_22/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4514 gnd OAI21X1_51/Y XNOR2X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4515 XNOR2X1_33/a_18_6# XNOR2X1_33/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4516 AOI22X1_48/D OAI21X1_51/Y XNOR2X1_33/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4517 XNOR2X1_33/a_35_6# XNOR2X1_33/a_2_6# AOI22X1_48/D Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4518 gnd AND2X2_22/Y XNOR2X1_33/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4519 XNOR2X1_33/a_12_41# AND2X2_22/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4520 AND2X2_22/a_2_6# XOR2X1_54/B vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4521 vdd XOR2X1_54/A AND2X2_22/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4522 AND2X2_22/Y AND2X2_22/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4523 AND2X2_22/a_9_6# XOR2X1_54/B AND2X2_22/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4524 gnd XOR2X1_54/A AND2X2_22/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4525 AND2X2_22/Y AND2X2_22/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4526 vdd XOR2X1_54/A XOR2X1_54/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4527 XOR2X1_54/a_18_54# XOR2X1_54/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4528 XOR2X1_54/Y XOR2X1_54/A XOR2X1_54/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4529 XOR2X1_54/a_35_54# XOR2X1_54/a_2_6# XOR2X1_54/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4530 vdd XOR2X1_54/B XOR2X1_54/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4531 XOR2X1_54/a_13_43# XOR2X1_54/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4532 gnd XOR2X1_54/A XOR2X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4533 XOR2X1_54/a_18_6# XOR2X1_54/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4534 XOR2X1_54/Y XOR2X1_54/a_2_6# XOR2X1_54/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4535 XOR2X1_54/a_35_6# XOR2X1_54/A XOR2X1_54/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4536 gnd XOR2X1_54/B XOR2X1_54/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4537 XOR2X1_54/a_13_43# XOR2X1_54/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4538 vdd INVX2_28/Y XOR2X1_53/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4539 XOR2X1_53/a_18_54# XOR2X1_53/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4540 XOR2X1_53/Y INVX2_28/Y XOR2X1_53/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4541 XOR2X1_53/a_35_54# XOR2X1_53/a_2_6# XOR2X1_53/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4542 vdd XOR2X1_17/B XOR2X1_53/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4543 XOR2X1_53/a_13_43# XOR2X1_17/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4544 gnd INVX2_28/Y XOR2X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4545 XOR2X1_53/a_18_6# XOR2X1_53/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4546 XOR2X1_53/Y XOR2X1_53/a_2_6# XOR2X1_53/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4547 XOR2X1_53/a_35_6# INVX2_28/Y XOR2X1_53/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4548 gnd XOR2X1_17/B XOR2X1_53/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4549 XOR2X1_53/a_13_43# XOR2X1_17/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4550 vdd XOR2X1_54/Y AOI22X1_49/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4551 AOI22X1_49/a_2_54# INVX2_92/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4552 AND2X2_21/B INVX2_94/Y AOI22X1_49/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4553 AOI22X1_49/a_2_54# XOR2X1_58/Y AND2X2_21/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4554 AOI22X1_49/a_11_6# XOR2X1_54/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4555 AND2X2_21/B INVX2_92/Y AOI22X1_49/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4556 AOI22X1_49/a_28_6# INVX2_94/Y AND2X2_21/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4557 gnd XOR2X1_58/Y AOI22X1_49/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4558 vdd INVX2_94/Y AOI22X1_48/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4559 AOI22X1_48/a_2_54# AOI22X1_48/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4560 AOI22X1_48/Y AOI22X1_48/D AOI22X1_48/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4561 AOI22X1_48/a_2_54# INVX2_92/Y AOI22X1_48/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4562 AOI22X1_48/a_11_6# INVX2_94/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4563 AOI22X1_48/Y AOI22X1_48/B AOI22X1_48/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4564 AOI22X1_48/a_28_6# AOI22X1_48/D AOI22X1_48/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4565 gnd INVX2_92/Y AOI22X1_48/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4566 AND2X2_21/a_2_6# AND2X2_21/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4567 vdd AND2X2_21/B AND2X2_21/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4568 AND2X2_21/Y AND2X2_21/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4569 AND2X2_21/a_9_6# AND2X2_21/A AND2X2_21/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4570 gnd AND2X2_21/B AND2X2_21/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4571 AND2X2_21/Y AND2X2_21/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4572 vdd OAI21X1_49/Y XNOR2X1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4573 XNOR2X1_30/a_18_54# XNOR2X1_30/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4574 AOI22X1_55/D XNOR2X1_30/a_2_6# XNOR2X1_30/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4575 XNOR2X1_30/a_35_54# OAI21X1_49/Y AOI22X1_55/D vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4576 vdd AND2X2_23/Y XNOR2X1_30/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4577 XNOR2X1_30/a_12_41# AND2X2_23/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4578 gnd OAI21X1_49/Y XNOR2X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4579 XNOR2X1_30/a_18_6# XNOR2X1_30/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4580 AOI22X1_55/D OAI21X1_49/Y XNOR2X1_30/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4581 XNOR2X1_30/a_35_6# XNOR2X1_30/a_2_6# AOI22X1_55/D Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4582 gnd AND2X2_23/Y XNOR2X1_30/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4583 XNOR2X1_30/a_12_41# AND2X2_23/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4584 OAI21X1_49/a_9_54# OAI21X1_56/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4585 OAI21X1_49/Y INVX2_67/Y OAI21X1_49/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4586 vdd NAND3X1_25/B OAI21X1_49/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4587 gnd OAI21X1_56/A OAI21X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4588 OAI21X1_49/a_2_6# INVX2_67/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4589 OAI21X1_49/Y NAND3X1_25/B OAI21X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4590 INVX2_67/Y INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4591 INVX2_67/Y INVX2_67/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4592 vdd BUFX2_11/Y DFFPOSX1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4593 DFFPOSX1_41/a_17_74# OAI22X1_8/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4594 DFFPOSX1_41/a_22_6# BUFX2_11/Y DFFPOSX1_41/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4595 DFFPOSX1_41/a_31_74# DFFPOSX1_41/a_2_6# DFFPOSX1_41/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4596 vdd DFFPOSX1_41/a_34_4# DFFPOSX1_41/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4597 DFFPOSX1_41/a_34_4# DFFPOSX1_41/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4598 DFFPOSX1_41/a_61_74# DFFPOSX1_41/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4599 DFFPOSX1_41/a_66_6# DFFPOSX1_41/a_2_6# DFFPOSX1_41/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4600 DFFPOSX1_41/a_76_84# BUFX2_11/Y DFFPOSX1_41/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4601 vdd INVX2_86/A DFFPOSX1_41/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4602 gnd BUFX2_11/Y DFFPOSX1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4603 INVX2_86/A DFFPOSX1_41/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4604 DFFPOSX1_41/a_17_6# OAI22X1_8/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4605 DFFPOSX1_41/a_22_6# DFFPOSX1_41/a_2_6# DFFPOSX1_41/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4606 DFFPOSX1_41/a_31_6# BUFX2_11/Y DFFPOSX1_41/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4607 gnd DFFPOSX1_41/a_34_4# DFFPOSX1_41/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4608 DFFPOSX1_41/a_34_4# DFFPOSX1_41/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4609 DFFPOSX1_41/a_61_6# DFFPOSX1_41/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4610 DFFPOSX1_41/a_66_6# BUFX2_11/Y DFFPOSX1_41/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4611 DFFPOSX1_41/a_76_6# DFFPOSX1_41/a_2_6# DFFPOSX1_41/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4612 gnd INVX2_86/A DFFPOSX1_41/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4613 INVX2_86/A DFFPOSX1_41/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4614 OAI22X1_8/a_9_54# INVX2_49/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4615 OAI22X1_8/Y INVX2_84/Y OAI22X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4616 OAI22X1_8/a_28_54# INVX2_99/Y OAI22X1_8/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4617 vdd INVX2_86/Y OAI22X1_8/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4618 gnd INVX2_49/Y OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4619 OAI22X1_8/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4620 OAI22X1_8/Y INVX2_99/Y OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4621 OAI22X1_8/a_2_6# INVX2_86/Y OAI22X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4622 OAI22X1_6/a_9_54# INVX2_63/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4623 OAI22X1_6/Y INVX2_84/Y OAI22X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4624 OAI22X1_6/a_28_54# INVX2_99/Y OAI22X1_6/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4625 vdd OAI22X1_6/C OAI22X1_6/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4626 gnd INVX2_63/Y OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4627 OAI22X1_6/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4628 OAI22X1_6/Y INVX2_99/Y OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4629 OAI22X1_6/a_2_6# OAI22X1_6/C OAI22X1_6/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4630 INVX2_66/Y INVX2_66/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4631 INVX2_66/Y INVX2_66/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4632 vdd INVX2_61/Y DFFPOSX1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4633 DFFPOSX1_38/a_17_74# INVX2_56/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4634 DFFPOSX1_38/a_22_6# INVX2_61/Y DFFPOSX1_38/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4635 DFFPOSX1_38/a_31_74# DFFPOSX1_38/a_2_6# DFFPOSX1_38/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4636 vdd DFFPOSX1_38/a_34_4# DFFPOSX1_38/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4637 DFFPOSX1_38/a_34_4# DFFPOSX1_38/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4638 DFFPOSX1_38/a_61_74# DFFPOSX1_38/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4639 DFFPOSX1_38/a_66_6# DFFPOSX1_38/a_2_6# DFFPOSX1_38/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4640 DFFPOSX1_38/a_76_84# INVX2_61/Y DFFPOSX1_38/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4641 vdd con_writeout DFFPOSX1_38/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4642 gnd INVX2_61/Y DFFPOSX1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4643 con_writeout DFFPOSX1_38/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4644 DFFPOSX1_38/a_17_6# INVX2_56/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4645 DFFPOSX1_38/a_22_6# DFFPOSX1_38/a_2_6# DFFPOSX1_38/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4646 DFFPOSX1_38/a_31_6# INVX2_61/Y DFFPOSX1_38/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4647 gnd DFFPOSX1_38/a_34_4# DFFPOSX1_38/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4648 DFFPOSX1_38/a_34_4# DFFPOSX1_38/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4649 DFFPOSX1_38/a_61_6# DFFPOSX1_38/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4650 DFFPOSX1_38/a_66_6# INVX2_61/Y DFFPOSX1_38/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4651 DFFPOSX1_38/a_76_6# DFFPOSX1_38/a_2_6# DFFPOSX1_38/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4652 gnd con_writeout DFFPOSX1_38/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4653 con_writeout DFFPOSX1_38/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4654 INVX2_63/Y INVX2_63/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4655 INVX2_63/Y INVX2_63/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4656 OAI22X1_4/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4657 OAI22X1_4/Y INVX2_63/Y OAI22X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4658 OAI22X1_4/a_28_54# INVX2_60/Y OAI22X1_4/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4659 vdd INVX2_62/Y OAI22X1_4/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4660 gnd BUFX2_3/Y OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4661 OAI22X1_4/a_2_6# INVX2_63/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4662 OAI22X1_4/Y INVX2_60/Y OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4663 OAI22X1_4/a_2_6# INVX2_62/Y OAI22X1_4/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4664 vdd BUFX2_8/A BUFX2_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4665 BUFX2_4/Y BUFX2_4/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4666 gnd BUFX2_8/A BUFX2_4/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4667 BUFX2_4/Y BUFX2_4/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4668 vdd BUFX2_8/A BUFX2_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4669 BUFX2_3/Y BUFX2_3/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4670 gnd BUFX2_8/A BUFX2_3/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4671 BUFX2_3/Y BUFX2_3/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4672 vdd BUFX2_8/A BUFX2_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4673 BUFX2_2/Y BUFX2_2/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4674 gnd BUFX2_8/A BUFX2_2/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M4675 BUFX2_2/Y BUFX2_2/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4676 INVX2_60/Y out_MemBData[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4677 INVX2_60/Y out_MemBData[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4678 vdd BUFX2_11/Y DFFPOSX1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4679 DFFPOSX1_36/a_17_74# OAI21X1_47/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4680 DFFPOSX1_36/a_22_6# BUFX2_11/Y DFFPOSX1_36/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4681 DFFPOSX1_36/a_31_74# DFFPOSX1_36/a_2_6# DFFPOSX1_36/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4682 vdd DFFPOSX1_36/a_34_4# DFFPOSX1_36/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4683 DFFPOSX1_36/a_34_4# DFFPOSX1_36/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4684 DFFPOSX1_36/a_61_74# DFFPOSX1_36/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4685 DFFPOSX1_36/a_66_6# DFFPOSX1_36/a_2_6# DFFPOSX1_36/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4686 DFFPOSX1_36/a_76_84# BUFX2_11/Y DFFPOSX1_36/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4687 vdd out_MemBData[2] DFFPOSX1_36/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4688 gnd BUFX2_11/Y DFFPOSX1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4689 out_MemBData[2] DFFPOSX1_36/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4690 DFFPOSX1_36/a_17_6# OAI21X1_47/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4691 DFFPOSX1_36/a_22_6# DFFPOSX1_36/a_2_6# DFFPOSX1_36/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4692 DFFPOSX1_36/a_31_6# BUFX2_11/Y DFFPOSX1_36/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4693 gnd DFFPOSX1_36/a_34_4# DFFPOSX1_36/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4694 DFFPOSX1_36/a_34_4# DFFPOSX1_36/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4695 DFFPOSX1_36/a_61_6# DFFPOSX1_36/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4696 DFFPOSX1_36/a_66_6# BUFX2_11/Y DFFPOSX1_36/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4697 DFFPOSX1_36/a_76_6# DFFPOSX1_36/a_2_6# DFFPOSX1_36/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4698 gnd out_MemBData[2] DFFPOSX1_36/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4699 out_MemBData[2] DFFPOSX1_36/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4700 AND2X2_19/a_2_6# OR2X2_0/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4701 vdd BUFX2_2/Y AND2X2_19/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4702 AND2X2_19/Y AND2X2_19/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4703 AND2X2_19/a_9_6# OR2X2_0/A AND2X2_19/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4704 gnd BUFX2_2/Y AND2X2_19/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4705 AND2X2_19/Y AND2X2_19/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4706 INVX2_58/Y con_readData vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4707 INVX2_58/Y con_readData gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4708 OAI21X1_46/a_9_54# INVX2_58/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4709 OAI21X1_45/B OAI21X1_46/B OAI21X1_46/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4710 vdd BUFX2_2/Y OAI21X1_45/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4711 gnd INVX2_58/Y OAI21X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4712 OAI21X1_46/a_2_6# OAI21X1_46/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4713 OAI21X1_45/B BUFX2_2/Y OAI21X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4714 OAI21X1_45/a_9_54# INVX2_57/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4715 OAI21X1_45/Y OAI21X1_45/B OAI21X1_45/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4716 vdd OAI21X1_45/C OAI21X1_45/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4717 gnd INVX2_57/Y OAI21X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4718 OAI21X1_45/a_2_6# OAI21X1_45/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4719 OAI21X1_45/Y OAI21X1_45/C OAI21X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4720 INVX2_57/Y INVX2_57/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4721 INVX2_57/Y INVX2_57/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4722 OAI21X1_43/a_9_54# con_readData vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4723 OR2X2_0/A con_loadData OAI21X1_43/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4724 vdd con_writeData OR2X2_0/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4725 gnd con_readData OAI21X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4726 OAI21X1_43/a_2_6# con_loadData gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4727 OR2X2_0/A con_writeData OAI21X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4728 OAI21X1_42/a_9_54# con_readData vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4729 INVX2_72/A con_loadData OAI21X1_42/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4730 vdd BUFX2_2/Y INVX2_72/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4731 gnd con_readData OAI21X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4732 OAI21X1_42/a_2_6# con_loadData gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4733 INVX2_72/A BUFX2_2/Y OAI21X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4734 INVX2_56/Y INVX2_56/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4735 INVX2_56/Y INVX2_56/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4736 vdd INVX2_43/Y DFFPOSX1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4737 DFFPOSX1_35/a_17_74# INVX2_55/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4738 DFFPOSX1_35/a_22_6# INVX2_43/Y DFFPOSX1_35/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4739 DFFPOSX1_35/a_31_74# DFFPOSX1_35/a_2_6# DFFPOSX1_35/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4740 vdd DFFPOSX1_35/a_34_4# DFFPOSX1_35/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4741 DFFPOSX1_35/a_34_4# DFFPOSX1_35/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4742 DFFPOSX1_35/a_61_74# DFFPOSX1_35/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4743 DFFPOSX1_35/a_66_6# DFFPOSX1_35/a_2_6# DFFPOSX1_35/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4744 DFFPOSX1_35/a_76_84# INVX2_43/Y DFFPOSX1_35/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4745 vdd con_loadData DFFPOSX1_35/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4746 gnd INVX2_43/Y DFFPOSX1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4747 con_loadData DFFPOSX1_35/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4748 DFFPOSX1_35/a_17_6# INVX2_55/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4749 DFFPOSX1_35/a_22_6# DFFPOSX1_35/a_2_6# DFFPOSX1_35/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4750 DFFPOSX1_35/a_31_6# INVX2_43/Y DFFPOSX1_35/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4751 gnd DFFPOSX1_35/a_34_4# DFFPOSX1_35/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4752 DFFPOSX1_35/a_34_4# DFFPOSX1_35/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4753 DFFPOSX1_35/a_61_6# DFFPOSX1_35/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4754 DFFPOSX1_35/a_66_6# INVX2_43/Y DFFPOSX1_35/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4755 DFFPOSX1_35/a_76_6# DFFPOSX1_35/a_2_6# DFFPOSX1_35/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4756 gnd con_loadData DFFPOSX1_35/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4757 con_loadData DFFPOSX1_35/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4758 INVX2_55/Y INVX2_55/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4759 INVX2_55/Y INVX2_55/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4760 INVX2_55/A INVX2_51/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4761 vdd INVX2_40/Y INVX2_55/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4762 INVX2_55/A INVX2_52/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4763 NAND3X1_19/a_9_6# INVX2_51/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4764 NAND3X1_19/a_14_6# INVX2_40/Y NAND3X1_19/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4765 INVX2_55/A INVX2_52/A NAND3X1_19/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4766 INVX2_52/Y INVX2_52/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4767 INVX2_52/Y INVX2_52/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4768 NAND3X1_22/B OAI21X1_50/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4769 vdd OAI21X1_50/B NAND3X1_22/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4770 NAND2X1_20/a_9_6# OAI21X1_50/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4771 NAND3X1_22/B OAI21X1_50/B NAND2X1_20/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4772 OAI21X1_51/a_9_54# OAI21X1_50/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4773 OAI21X1_51/Y OAI21X1_50/B OAI21X1_51/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4774 vdd NAND3X1_22/B OAI21X1_51/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4775 gnd OAI21X1_50/A OAI21X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4776 OAI21X1_51/a_2_6# OAI21X1_50/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4777 OAI21X1_51/Y NAND3X1_22/B OAI21X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4778 OAI21X1_50/a_9_54# OAI21X1_50/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4779 XOR2X1_49/A OAI21X1_50/B OAI21X1_50/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4780 vdd NAND3X1_22/Y XOR2X1_49/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4781 gnd OAI21X1_50/A OAI21X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4782 OAI21X1_50/a_2_6# OAI21X1_50/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4783 XOR2X1_49/A NAND3X1_22/Y OAI21X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4784 NAND3X1_22/Y XOR2X1_54/B vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4785 vdd NAND3X1_22/B NAND3X1_22/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4786 NAND3X1_22/Y XOR2X1_54/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4787 NAND3X1_22/a_9_6# XOR2X1_54/B gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4788 NAND3X1_22/a_14_6# NAND3X1_22/B NAND3X1_22/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4789 NAND3X1_22/Y XOR2X1_54/A NAND3X1_22/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4790 vdd XOR2X1_17/B XNOR2X1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4791 XNOR2X1_32/a_18_54# XNOR2X1_32/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4792 XOR2X1_54/B XNOR2X1_32/a_2_6# XNOR2X1_32/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4793 XNOR2X1_32/a_35_54# XOR2X1_17/B XOR2X1_54/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4794 vdd XOR2X1_48/Y XNOR2X1_32/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4795 XNOR2X1_32/a_12_41# XOR2X1_48/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4796 gnd XOR2X1_17/B XNOR2X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4797 XNOR2X1_32/a_18_6# XNOR2X1_32/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4798 XOR2X1_54/B XOR2X1_17/B XNOR2X1_32/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4799 XNOR2X1_32/a_35_6# XNOR2X1_32/a_2_6# XOR2X1_54/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4800 gnd XOR2X1_48/Y XNOR2X1_32/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4801 XNOR2X1_32/a_12_41# XOR2X1_48/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4802 vdd XOR2X1_81/A XNOR2X1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4803 XNOR2X1_31/a_18_54# XNOR2X1_31/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4804 XOR2X1_54/A XNOR2X1_31/a_2_6# XNOR2X1_31/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4805 XNOR2X1_31/a_35_54# XOR2X1_81/A XOR2X1_54/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4806 vdd XOR2X1_51/Y XNOR2X1_31/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4807 XNOR2X1_31/a_12_41# XOR2X1_51/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4808 gnd XOR2X1_81/A XNOR2X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4809 XNOR2X1_31/a_18_6# XNOR2X1_31/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4810 XOR2X1_54/A XOR2X1_81/A XNOR2X1_31/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4811 XNOR2X1_31/a_35_6# XNOR2X1_31/a_2_6# XOR2X1_54/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4812 gnd XOR2X1_51/Y XNOR2X1_31/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4813 XNOR2X1_31/a_12_41# XOR2X1_51/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4814 vdd out_MuxData[11] AOI22X1_47/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M4815 AOI22X1_47/a_2_54# out_MuxData[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4816 OAI21X1_50/A out_MuxData[1] AOI22X1_47/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M4817 AOI22X1_47/a_2_54# XOR2X1_51/Y OAI21X1_50/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4818 AOI22X1_47/a_11_6# out_MuxData[11] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4819 OAI21X1_50/A out_MuxData[13] AOI22X1_47/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4820 AOI22X1_47/a_28_6# out_MuxData[1] OAI21X1_50/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4821 gnd XOR2X1_51/Y AOI22X1_47/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4822 vdd OAI22X1_6/C XOR2X1_52/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4823 XOR2X1_52/a_18_54# XOR2X1_52/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4824 XOR2X1_52/Y OAI22X1_6/C XOR2X1_52/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4825 XOR2X1_52/a_35_54# XOR2X1_52/a_2_6# XOR2X1_52/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4826 vdd INVX2_86/Y XOR2X1_52/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4827 XOR2X1_52/a_13_43# INVX2_86/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4828 gnd OAI22X1_6/C XOR2X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4829 XOR2X1_52/a_18_6# XOR2X1_52/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4830 XOR2X1_52/Y XOR2X1_52/a_2_6# XOR2X1_52/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4831 XOR2X1_52/a_35_6# OAI22X1_6/C XOR2X1_52/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4832 gnd INVX2_86/Y XOR2X1_52/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4833 XOR2X1_52/a_13_43# INVX2_86/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4834 vdd INVX2_50/Y XOR2X1_51/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4835 XOR2X1_51/a_18_54# XOR2X1_51/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4836 XOR2X1_51/Y INVX2_50/Y XOR2X1_51/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4837 XOR2X1_51/a_35_54# XOR2X1_51/a_2_6# XOR2X1_51/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4838 vdd INVX2_87/Y XOR2X1_51/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4839 XOR2X1_51/a_13_43# INVX2_87/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4840 gnd INVX2_50/Y XOR2X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4841 XOR2X1_51/a_18_6# XOR2X1_51/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4842 XOR2X1_51/Y XOR2X1_51/a_2_6# XOR2X1_51/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4843 XOR2X1_51/a_35_6# INVX2_50/Y XOR2X1_51/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4844 gnd INVX2_87/Y XOR2X1_51/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4845 XOR2X1_51/a_13_43# INVX2_87/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4846 NOR2X1_16/A AOI22X1_48/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M4847 vdd AOI22X1_55/Y NOR2X1_16/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4848 NOR2X1_16/A AND2X2_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4849 NAND3X1_21/a_9_6# AOI22X1_48/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4850 NAND3X1_21/a_14_6# AOI22X1_55/Y NAND3X1_21/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M4851 NOR2X1_16/A AND2X2_13/Y NAND3X1_21/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M4852 vdd INVX2_86/Y XNOR2X1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4853 XNOR2X1_29/a_18_54# XNOR2X1_29/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4854 XOR2X1_55/A XNOR2X1_29/a_2_6# XNOR2X1_29/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M4855 XNOR2X1_29/a_35_54# INVX2_86/Y XOR2X1_55/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4856 vdd XOR2X1_46/Y XNOR2X1_29/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4857 XNOR2X1_29/a_12_41# XOR2X1_46/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4858 gnd INVX2_86/Y XNOR2X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4859 XNOR2X1_29/a_18_6# XNOR2X1_29/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4860 XOR2X1_55/A INVX2_86/Y XNOR2X1_29/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M4861 XNOR2X1_29/a_35_6# XNOR2X1_29/a_2_6# XOR2X1_55/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4862 gnd XOR2X1_46/Y XNOR2X1_29/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4863 XNOR2X1_29/a_12_41# XOR2X1_46/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4864 NAND3X1_25/B OAI21X1_56/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4865 vdd INVX2_67/Y NAND3X1_25/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4866 NAND2X1_19/a_9_6# OAI21X1_56/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4867 NAND3X1_25/B INVX2_67/Y NAND2X1_19/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4868 AND2X2_20/a_2_6# AND2X2_20/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4869 vdd AND2X2_20/B AND2X2_20/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4870 AND2X2_20/Y AND2X2_20/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4871 AND2X2_20/a_9_6# AND2X2_20/A AND2X2_20/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M4872 gnd AND2X2_20/B AND2X2_20/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4873 AND2X2_20/Y AND2X2_20/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4874 vdd BUFX2_11/Y DFFPOSX1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4875 DFFPOSX1_40/a_17_74# OAI22X1_7/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4876 DFFPOSX1_40/a_22_6# BUFX2_11/Y DFFPOSX1_40/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4877 DFFPOSX1_40/a_31_74# DFFPOSX1_40/a_2_6# DFFPOSX1_40/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4878 vdd DFFPOSX1_40/a_34_4# DFFPOSX1_40/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4879 DFFPOSX1_40/a_34_4# DFFPOSX1_40/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4880 DFFPOSX1_40/a_61_74# DFFPOSX1_40/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4881 DFFPOSX1_40/a_66_6# DFFPOSX1_40/a_2_6# DFFPOSX1_40/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4882 DFFPOSX1_40/a_76_84# BUFX2_11/Y DFFPOSX1_40/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4883 vdd out_MuxData[1] DFFPOSX1_40/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4884 gnd BUFX2_11/Y DFFPOSX1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4885 out_MuxData[1] DFFPOSX1_40/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4886 DFFPOSX1_40/a_17_6# OAI22X1_7/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4887 DFFPOSX1_40/a_22_6# DFFPOSX1_40/a_2_6# DFFPOSX1_40/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4888 DFFPOSX1_40/a_31_6# BUFX2_11/Y DFFPOSX1_40/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4889 gnd DFFPOSX1_40/a_34_4# DFFPOSX1_40/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4890 DFFPOSX1_40/a_34_4# DFFPOSX1_40/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4891 DFFPOSX1_40/a_61_6# DFFPOSX1_40/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4892 DFFPOSX1_40/a_66_6# BUFX2_11/Y DFFPOSX1_40/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4893 DFFPOSX1_40/a_76_6# DFFPOSX1_40/a_2_6# DFFPOSX1_40/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4894 gnd out_MuxData[1] DFFPOSX1_40/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4895 out_MuxData[1] DFFPOSX1_40/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4896 OAI22X1_7/a_9_54# INVX2_48/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4897 OAI22X1_7/Y INVX2_84/Y OAI22X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4898 OAI22X1_7/a_28_54# INVX2_99/Y OAI22X1_7/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4899 vdd XOR2X1_81/A OAI22X1_7/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4900 gnd INVX2_48/Y OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4901 OAI22X1_7/a_2_6# INVX2_84/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4902 OAI22X1_7/Y INVX2_99/Y OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4903 OAI22X1_7/a_2_6# XOR2X1_81/A OAI22X1_7/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4904 vdd BUFX2_5/Y DFFPOSX1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4905 DFFPOSX1_39/a_17_74# INVX2_66/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4906 DFFPOSX1_39/a_22_6# BUFX2_5/Y DFFPOSX1_39/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4907 DFFPOSX1_39/a_31_74# DFFPOSX1_39/a_2_6# DFFPOSX1_39/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4908 vdd DFFPOSX1_39/a_34_4# DFFPOSX1_39/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4909 DFFPOSX1_39/a_34_4# DFFPOSX1_39/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4910 DFFPOSX1_39/a_61_74# DFFPOSX1_39/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4911 DFFPOSX1_39/a_66_6# DFFPOSX1_39/a_2_6# DFFPOSX1_39/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4912 DFFPOSX1_39/a_76_84# BUFX2_5/Y DFFPOSX1_39/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4913 vdd INVX2_39/A DFFPOSX1_39/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4914 gnd BUFX2_5/Y DFFPOSX1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4915 INVX2_39/A DFFPOSX1_39/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4916 DFFPOSX1_39/a_17_6# INVX2_66/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4917 DFFPOSX1_39/a_22_6# DFFPOSX1_39/a_2_6# DFFPOSX1_39/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4918 DFFPOSX1_39/a_31_6# BUFX2_5/Y DFFPOSX1_39/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4919 gnd DFFPOSX1_39/a_34_4# DFFPOSX1_39/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4920 DFFPOSX1_39/a_34_4# DFFPOSX1_39/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4921 DFFPOSX1_39/a_61_6# DFFPOSX1_39/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4922 DFFPOSX1_39/a_66_6# BUFX2_5/Y DFFPOSX1_39/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4923 DFFPOSX1_39/a_76_6# DFFPOSX1_39/a_2_6# DFFPOSX1_39/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4924 gnd INVX2_39/A DFFPOSX1_39/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4925 INVX2_39/A DFFPOSX1_39/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4926 INVX2_65/Y INVX2_65/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4927 INVX2_65/Y INVX2_65/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4928 OAI22X1_5/a_9_54# BUFX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4929 OAI22X1_5/Y INVX2_65/Y OAI22X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4930 OAI22X1_5/a_28_54# INVX2_64/Y OAI22X1_5/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4931 vdd INVX2_62/Y OAI22X1_5/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4932 gnd BUFX2_4/Y OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4933 OAI22X1_5/a_2_6# INVX2_65/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4934 OAI22X1_5/Y INVX2_64/Y OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4935 OAI22X1_5/a_2_6# INVX2_62/Y OAI22X1_5/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4936 INVX2_64/Y out_MemBData[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4937 INVX2_64/Y out_MemBData[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4938 vdd in_clkb DFFPOSX1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M4939 DFFPOSX1_37/a_17_74# OAI22X1_4/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4940 DFFPOSX1_37/a_22_6# in_clkb DFFPOSX1_37/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4941 DFFPOSX1_37/a_31_74# DFFPOSX1_37/a_2_6# DFFPOSX1_37/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M4942 vdd DFFPOSX1_37/a_34_4# DFFPOSX1_37/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4943 DFFPOSX1_37/a_34_4# DFFPOSX1_37/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4944 DFFPOSX1_37/a_61_74# DFFPOSX1_37/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4945 DFFPOSX1_37/a_66_6# DFFPOSX1_37/a_2_6# DFFPOSX1_37/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M4946 DFFPOSX1_37/a_76_84# in_clkb DFFPOSX1_37/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4947 vdd INVX2_63/A DFFPOSX1_37/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4948 gnd in_clkb DFFPOSX1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M4949 INVX2_63/A DFFPOSX1_37/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4950 DFFPOSX1_37/a_17_6# OAI22X1_4/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4951 DFFPOSX1_37/a_22_6# DFFPOSX1_37/a_2_6# DFFPOSX1_37/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4952 DFFPOSX1_37/a_31_6# in_clkb DFFPOSX1_37/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4953 gnd DFFPOSX1_37/a_34_4# DFFPOSX1_37/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4954 DFFPOSX1_37/a_34_4# DFFPOSX1_37/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M4955 DFFPOSX1_37/a_61_6# DFFPOSX1_37/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4956 DFFPOSX1_37/a_66_6# in_clkb DFFPOSX1_37/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M4957 DFFPOSX1_37/a_76_6# DFFPOSX1_37/a_2_6# DFFPOSX1_37/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M4958 gnd INVX2_63/A DFFPOSX1_37/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4959 INVX2_63/A DFFPOSX1_37/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4960 INVX2_62/Y BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4961 INVX2_62/Y BUFX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4962 INVX2_61/Y BUFX2_1/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4963 INVX2_61/Y BUFX2_1/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4964 OAI21X1_48/a_9_54# NOR2X1_13/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4965 OAI21X1_47/C AND2X2_19/Y OAI21X1_48/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4966 vdd out_MemBData[2] OAI21X1_47/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4967 gnd NOR2X1_13/Y OAI21X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4968 OAI21X1_48/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4969 OAI21X1_47/C out_MemBData[2] OAI21X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4970 OAI21X1_47/a_9_54# INVX2_59/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4971 OAI21X1_47/Y OR2X2_0/Y OAI21X1_47/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4972 vdd OAI21X1_47/C OAI21X1_47/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4973 gnd INVX2_59/A OAI21X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M4974 OAI21X1_47/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4975 OAI21X1_47/Y OAI21X1_47/C OAI21X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4976 INVX2_59/Y INVX2_59/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4977 INVX2_59/Y INVX2_59/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4978 OR2X2_0/a_9_54# OR2X2_0/A OR2X2_0/a_2_54# vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M4979 vdd OR2X2_0/B OR2X2_0/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4980 OR2X2_0/Y OR2X2_0/a_2_54# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M4981 OR2X2_0/a_2_54# OR2X2_0/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M4982 gnd OR2X2_0/B OR2X2_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4983 OR2X2_0/Y OR2X2_0/a_2_54# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4984 OAI21X1_46/B con_writeData vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4985 vdd INVX2_71/Y OAI21X1_46/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4986 NAND2X1_18/a_9_6# con_writeData gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M4987 OAI21X1_46/B INVX2_71/Y NAND2X1_18/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M4988 OAI22X1_3/a_9_54# con_readData vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4989 OR2X2_0/B in_DataIn OAI22X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M4990 OAI22X1_3/a_28_54# INVX2_58/Y OR2X2_0/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4991 vdd OAI22X1_3/C OAI22X1_3/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4992 gnd con_readData OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M4993 OAI22X1_3/a_2_6# in_DataIn gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4994 OR2X2_0/B INVX2_58/Y OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M4995 OAI22X1_3/a_2_6# OAI22X1_3/C OR2X2_0/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4996 OAI21X1_44/a_9_54# con_readData vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M4997 NAND2X1_17/B INVX2_54/Y OAI21X1_44/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M4998 vdd OAI21X1_44/C NAND2X1_17/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4999 gnd con_readData OAI21X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5000 OAI21X1_44/a_2_6# INVX2_54/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5001 NAND2X1_17/B OAI21X1_44/C OAI21X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5002 OAI21X1_45/C con_writeData vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5003 vdd NAND2X1_17/B OAI21X1_45/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5004 NAND2X1_17/a_9_6# con_writeData gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5005 OAI21X1_45/C NAND2X1_17/B NAND2X1_17/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5006 INVX2_54/Y con_loadData vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5007 INVX2_54/Y con_loadData gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5008 vdd INVX2_43/Y DFFPOSX1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5009 DFFPOSX1_34/a_17_74# INVX2_53/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5010 DFFPOSX1_34/a_22_6# INVX2_43/Y DFFPOSX1_34/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5011 DFFPOSX1_34/a_31_74# DFFPOSX1_34/a_2_6# DFFPOSX1_34/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5012 vdd DFFPOSX1_34/a_34_4# DFFPOSX1_34/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5013 DFFPOSX1_34/a_34_4# DFFPOSX1_34/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5014 DFFPOSX1_34/a_61_74# DFFPOSX1_34/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5015 DFFPOSX1_34/a_66_6# DFFPOSX1_34/a_2_6# DFFPOSX1_34/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5016 DFFPOSX1_34/a_76_84# INVX2_43/Y DFFPOSX1_34/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5017 vdd con_writeData DFFPOSX1_34/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5018 gnd INVX2_43/Y DFFPOSX1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5019 con_writeData DFFPOSX1_34/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5020 DFFPOSX1_34/a_17_6# INVX2_53/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5021 DFFPOSX1_34/a_22_6# DFFPOSX1_34/a_2_6# DFFPOSX1_34/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5022 DFFPOSX1_34/a_31_6# INVX2_43/Y DFFPOSX1_34/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5023 gnd DFFPOSX1_34/a_34_4# DFFPOSX1_34/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5024 DFFPOSX1_34/a_34_4# DFFPOSX1_34/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5025 DFFPOSX1_34/a_61_6# DFFPOSX1_34/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5026 DFFPOSX1_34/a_66_6# INVX2_43/Y DFFPOSX1_34/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5027 DFFPOSX1_34/a_76_6# DFFPOSX1_34/a_2_6# DFFPOSX1_34/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5028 gnd con_writeData DFFPOSX1_34/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5029 con_writeData DFFPOSX1_34/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5030 INVX2_53/Y INVX2_53/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5031 INVX2_53/Y INVX2_53/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5032 INVX2_11/A INVX2_56/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5033 vdd OAI21X1_52/C INVX2_11/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5034 NAND2X1_16/a_9_6# INVX2_56/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5035 INVX2_11/A OAI21X1_52/C NAND2X1_16/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5036 OAI21X1_52/C INVX2_52/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5037 vdd INVX2_51/A OAI21X1_52/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5038 OAI21X1_52/C INVX2_40/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5039 NAND3X1_20/a_9_6# INVX2_52/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5040 NAND3X1_20/a_14_6# INVX2_51/A NAND3X1_20/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5041 OAI21X1_52/C INVX2_40/A NAND3X1_20/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5042 INVX2_56/A INVX2_51/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5043 vdd INVX2_52/Y INVX2_56/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5044 INVX2_56/A INVX2_40/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5045 NAND3X1_18/a_9_6# INVX2_51/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5046 NAND3X1_18/a_14_6# INVX2_52/Y NAND3X1_18/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5047 INVX2_56/A INVX2_40/A NAND3X1_18/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5048 INVX2_51/Y INVX2_51/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5049 INVX2_51/Y INVX2_51/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5050 vdd NOR2X1_17/B XNOR2X1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5051 XNOR2X1_28/a_18_54# XNOR2X1_28/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5052 OAI21X1_50/B XNOR2X1_28/a_2_6# XNOR2X1_28/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5053 XNOR2X1_28/a_35_54# NOR2X1_17/B OAI21X1_50/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5054 vdd NOR2X1_17/A XNOR2X1_28/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5055 XNOR2X1_28/a_12_41# NOR2X1_17/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5056 gnd NOR2X1_17/B XNOR2X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5057 XNOR2X1_28/a_18_6# XNOR2X1_28/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5058 OAI21X1_50/B NOR2X1_17/B XNOR2X1_28/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5059 XNOR2X1_28/a_35_6# XNOR2X1_28/a_2_6# OAI21X1_50/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5060 gnd NOR2X1_17/A XNOR2X1_28/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5061 XNOR2X1_28/a_12_41# NOR2X1_17/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5062 vdd XOR2X1_49/A XOR2X1_49/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5063 XOR2X1_49/a_18_54# XOR2X1_49/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5064 XOR2X1_49/Y XOR2X1_49/A XOR2X1_49/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5065 XOR2X1_49/a_35_54# XOR2X1_49/a_2_6# XOR2X1_49/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5066 vdd NOR2X1_17/Y XOR2X1_49/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5067 XOR2X1_49/a_13_43# NOR2X1_17/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5068 gnd XOR2X1_49/A XOR2X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5069 XOR2X1_49/a_18_6# XOR2X1_49/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5070 XOR2X1_49/Y XOR2X1_49/a_2_6# XOR2X1_49/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5071 XOR2X1_49/a_35_6# XOR2X1_49/A XOR2X1_49/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5072 gnd NOR2X1_17/Y XOR2X1_49/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5073 XOR2X1_49/a_13_43# NOR2X1_17/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5074 vdd XOR2X1_48/B AOI22X1_46/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5075 AOI22X1_46/a_2_54# out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5076 NOR2X1_17/A out_MuxData[8] AOI22X1_46/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5077 AOI22X1_46/a_2_54# XOR2X1_48/Y NOR2X1_17/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5078 AOI22X1_46/a_11_6# XOR2X1_48/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5079 NOR2X1_17/A out_MuxData[9] AOI22X1_46/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5080 AOI22X1_46/a_28_6# out_MuxData[8] NOR2X1_17/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5081 gnd XOR2X1_48/Y AOI22X1_46/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5082 vdd out_MuxData[9] XOR2X1_48/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5083 XOR2X1_48/a_18_54# XOR2X1_48/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5084 XOR2X1_48/Y out_MuxData[9] XOR2X1_48/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5085 XOR2X1_48/a_35_54# XOR2X1_48/a_2_6# XOR2X1_48/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5086 vdd XOR2X1_48/B XOR2X1_48/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5087 XOR2X1_48/a_13_43# XOR2X1_48/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5088 gnd out_MuxData[9] XOR2X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5089 XOR2X1_48/a_18_6# XOR2X1_48/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5090 XOR2X1_48/Y XOR2X1_48/a_2_6# XOR2X1_48/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5091 XOR2X1_48/a_35_6# out_MuxData[9] XOR2X1_48/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5092 gnd XOR2X1_48/B XOR2X1_48/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5093 XOR2X1_48/a_13_43# XOR2X1_48/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5094 vdd out_MuxData[0] AOI22X1_45/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5095 AOI22X1_45/a_2_54# out_MuxData[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5096 NOR2X1_17/B out_MuxData[15] AOI22X1_45/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5097 AOI22X1_45/a_2_54# XOR2X1_52/Y NOR2X1_17/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5098 AOI22X1_45/a_11_6# out_MuxData[0] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5099 NOR2X1_17/B out_MuxData[3] AOI22X1_45/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5100 AOI22X1_45/a_28_6# out_MuxData[15] NOR2X1_17/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5101 gnd XOR2X1_52/Y AOI22X1_45/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5102 vdd INVX2_50/Y XOR2X1_47/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5103 XOR2X1_47/a_18_54# XOR2X1_47/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5104 XOR2X1_47/Y INVX2_50/Y XOR2X1_47/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5105 XOR2X1_47/a_35_54# XOR2X1_47/a_2_6# XOR2X1_47/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5106 vdd INVX2_86/Y XOR2X1_47/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5107 XOR2X1_47/a_13_43# INVX2_86/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5108 gnd INVX2_50/Y XOR2X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5109 XOR2X1_47/a_18_6# XOR2X1_47/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5110 XOR2X1_47/Y XOR2X1_47/a_2_6# XOR2X1_47/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5111 XOR2X1_47/a_35_6# INVX2_50/Y XOR2X1_47/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5112 gnd INVX2_86/Y XOR2X1_47/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5113 XOR2X1_47/a_13_43# INVX2_86/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5114 vdd INVX2_59/Y AOI22X1_44/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5115 AOI22X1_44/a_2_54# XOR2X1_50/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5116 AOI22X1_44/Y XOR2X1_57/Y AOI22X1_44/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5117 AOI22X1_44/a_2_54# INVX2_73/Y AOI22X1_44/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5118 AOI22X1_44/a_11_6# INVX2_59/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5119 AOI22X1_44/Y XOR2X1_50/Y AOI22X1_44/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5120 AOI22X1_44/a_28_6# XOR2X1_57/Y AOI22X1_44/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5121 gnd INVX2_73/Y AOI22X1_44/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5122 NOR2X1_16/a_9_54# NOR2X1_16/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5123 INVX2_46/A NOR2X1_16/B NOR2X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5124 INVX2_46/A NOR2X1_16/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5125 gnd NOR2X1_16/B INVX2_46/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5126 vdd out_MuxData[9] AOI22X1_43/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5127 AOI22X1_43/a_2_54# out_MuxData[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5128 OAI21X1_56/A out_MuxData[3] AOI22X1_43/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5129 AOI22X1_43/a_2_54# XOR2X1_46/Y OAI21X1_56/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5130 AOI22X1_43/a_11_6# out_MuxData[9] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5131 OAI21X1_56/A out_MuxData[15] AOI22X1_43/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5132 AOI22X1_43/a_28_6# out_MuxData[3] OAI21X1_56/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5133 gnd XOR2X1_46/Y AOI22X1_43/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5134 vdd XOR2X1_2/Y AOI22X1_42/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5135 AOI22X1_42/a_2_54# INVX2_93/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5136 AND2X2_20/B INVX2_92/Y AOI22X1_42/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5137 AOI22X1_42/a_2_54# XOR2X1_49/Y AND2X2_20/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5138 AOI22X1_42/a_11_6# XOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5139 AND2X2_20/B INVX2_93/Y AOI22X1_42/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5140 AOI22X1_42/a_28_6# INVX2_92/Y AND2X2_20/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5141 gnd XOR2X1_49/Y AOI22X1_42/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5142 vdd INVX2_87/Y XNOR2X1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5143 XNOR2X1_25/a_18_54# XNOR2X1_25/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5144 XOR2X1_37/B XNOR2X1_25/a_2_6# XNOR2X1_25/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5145 XNOR2X1_25/a_35_54# INVX2_87/Y XOR2X1_37/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5146 vdd XOR2X1_45/Y XNOR2X1_25/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5147 XNOR2X1_25/a_12_41# XOR2X1_45/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5148 gnd INVX2_87/Y XNOR2X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5149 XNOR2X1_25/a_18_6# XNOR2X1_25/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5150 XOR2X1_37/B INVX2_87/Y XNOR2X1_25/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5151 XNOR2X1_25/a_35_6# XNOR2X1_25/a_2_6# XOR2X1_37/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5152 gnd XOR2X1_45/Y XNOR2X1_25/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5153 XNOR2X1_25/a_12_41# XOR2X1_45/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5154 vdd out_MuxData[12] XOR2X1_45/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5155 XOR2X1_45/a_18_54# XOR2X1_45/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5156 XOR2X1_45/Y out_MuxData[12] XOR2X1_45/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5157 XOR2X1_45/a_35_54# XOR2X1_45/a_2_6# XOR2X1_45/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5158 vdd INVX2_39/A XOR2X1_45/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5159 XOR2X1_45/a_13_43# INVX2_39/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5160 gnd out_MuxData[12] XOR2X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5161 XOR2X1_45/a_18_6# XOR2X1_45/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5162 XOR2X1_45/Y XOR2X1_45/a_2_6# XOR2X1_45/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5163 XOR2X1_45/a_35_6# out_MuxData[12] XOR2X1_45/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5164 gnd INVX2_39/A XOR2X1_45/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5165 XOR2X1_45/a_13_43# INVX2_39/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5166 vdd out_MuxData[12] AOI22X1_39/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5167 AOI22X1_39/a_2_54# out_MuxData[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5168 NOR2X1_14/B out_MuxData[11] AOI22X1_39/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5169 AOI22X1_39/a_2_54# XOR2X1_45/Y NOR2X1_14/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5170 AOI22X1_39/a_11_6# out_MuxData[12] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5171 NOR2X1_14/B out_MuxData[15] AOI22X1_39/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5172 AOI22X1_39/a_28_6# out_MuxData[11] NOR2X1_14/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5173 gnd XOR2X1_45/Y AOI22X1_39/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5174 NOR2X1_14/a_9_54# NOR2X1_14/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5175 NOR2X1_14/Y NOR2X1_14/B NOR2X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5176 NOR2X1_14/Y NOR2X1_14/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5177 gnd NOR2X1_14/B NOR2X1_14/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5178 vdd in_clkb DFFPOSX1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5179 DFFPOSX1_33/a_17_74# OAI22X1_5/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5180 DFFPOSX1_33/a_22_6# in_clkb DFFPOSX1_33/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5181 DFFPOSX1_33/a_31_74# DFFPOSX1_33/a_2_6# DFFPOSX1_33/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5182 vdd DFFPOSX1_33/a_34_4# DFFPOSX1_33/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5183 DFFPOSX1_33/a_34_4# DFFPOSX1_33/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5184 DFFPOSX1_33/a_61_74# DFFPOSX1_33/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5185 DFFPOSX1_33/a_66_6# DFFPOSX1_33/a_2_6# DFFPOSX1_33/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5186 DFFPOSX1_33/a_76_84# in_clkb DFFPOSX1_33/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5187 vdd INVX2_65/A DFFPOSX1_33/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5188 gnd in_clkb DFFPOSX1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5189 INVX2_65/A DFFPOSX1_33/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5190 DFFPOSX1_33/a_17_6# OAI22X1_5/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5191 DFFPOSX1_33/a_22_6# DFFPOSX1_33/a_2_6# DFFPOSX1_33/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5192 DFFPOSX1_33/a_31_6# in_clkb DFFPOSX1_33/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5193 gnd DFFPOSX1_33/a_34_4# DFFPOSX1_33/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5194 DFFPOSX1_33/a_34_4# DFFPOSX1_33/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5195 DFFPOSX1_33/a_61_6# DFFPOSX1_33/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5196 DFFPOSX1_33/a_66_6# in_clkb DFFPOSX1_33/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5197 DFFPOSX1_33/a_76_6# DFFPOSX1_33/a_2_6# DFFPOSX1_33/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5198 gnd INVX2_65/A DFFPOSX1_33/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5199 INVX2_65/A DFFPOSX1_33/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5200 INVX2_49/Y INVX2_49/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5201 INVX2_49/Y INVX2_49/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5202 vdd in_clkb DFFPOSX1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5203 DFFPOSX1_31/a_17_74# OAI22X1_2/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5204 DFFPOSX1_31/a_22_6# in_clkb DFFPOSX1_31/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5205 DFFPOSX1_31/a_31_74# DFFPOSX1_31/a_2_6# DFFPOSX1_31/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5206 vdd DFFPOSX1_31/a_34_4# DFFPOSX1_31/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5207 DFFPOSX1_31/a_34_4# DFFPOSX1_31/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5208 DFFPOSX1_31/a_61_74# DFFPOSX1_31/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5209 DFFPOSX1_31/a_66_6# DFFPOSX1_31/a_2_6# DFFPOSX1_31/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5210 DFFPOSX1_31/a_76_84# in_clkb DFFPOSX1_31/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5211 vdd INVX2_49/A DFFPOSX1_31/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5212 gnd in_clkb DFFPOSX1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5213 INVX2_49/A DFFPOSX1_31/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5214 DFFPOSX1_31/a_17_6# OAI22X1_2/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5215 DFFPOSX1_31/a_22_6# DFFPOSX1_31/a_2_6# DFFPOSX1_31/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5216 DFFPOSX1_31/a_31_6# in_clkb DFFPOSX1_31/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5217 gnd DFFPOSX1_31/a_34_4# DFFPOSX1_31/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5218 DFFPOSX1_31/a_34_4# DFFPOSX1_31/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5219 DFFPOSX1_31/a_61_6# DFFPOSX1_31/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5220 DFFPOSX1_31/a_66_6# in_clkb DFFPOSX1_31/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5221 DFFPOSX1_31/a_76_6# DFFPOSX1_31/a_2_6# DFFPOSX1_31/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5222 gnd INVX2_49/A DFFPOSX1_31/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5223 INVX2_49/A DFFPOSX1_31/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5224 OAI22X1_2/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5225 OAI22X1_2/Y INVX2_49/Y OAI22X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M5226 OAI22X1_2/a_28_54# INVX2_38/Y OAI22X1_2/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5227 vdd INVX2_62/Y OAI22X1_2/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5228 gnd BUFX2_3/Y OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M5229 OAI22X1_2/a_2_6# INVX2_49/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5230 OAI22X1_2/Y INVX2_38/Y OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5231 OAI22X1_2/a_2_6# INVX2_62/Y OAI22X1_2/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5232 vdd in_clkb DFFPOSX1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5233 DFFPOSX1_30/a_17_74# OAI21X1_39/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5234 DFFPOSX1_30/a_22_6# in_clkb DFFPOSX1_30/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5235 DFFPOSX1_30/a_31_74# DFFPOSX1_30/a_2_6# DFFPOSX1_30/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5236 vdd DFFPOSX1_30/a_34_4# DFFPOSX1_30/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5237 DFFPOSX1_30/a_34_4# DFFPOSX1_30/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5238 DFFPOSX1_30/a_61_74# DFFPOSX1_30/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5239 DFFPOSX1_30/a_66_6# DFFPOSX1_30/a_2_6# DFFPOSX1_30/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5240 DFFPOSX1_30/a_76_84# in_clkb DFFPOSX1_30/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5241 vdd out_temp_addNum[0] DFFPOSX1_30/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5242 gnd in_clkb DFFPOSX1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5243 out_temp_addNum[0] DFFPOSX1_30/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5244 DFFPOSX1_30/a_17_6# OAI21X1_39/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5245 DFFPOSX1_30/a_22_6# DFFPOSX1_30/a_2_6# DFFPOSX1_30/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5246 DFFPOSX1_30/a_31_6# in_clkb DFFPOSX1_30/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5247 gnd DFFPOSX1_30/a_34_4# DFFPOSX1_30/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5248 DFFPOSX1_30/a_34_4# DFFPOSX1_30/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5249 DFFPOSX1_30/a_61_6# DFFPOSX1_30/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5250 DFFPOSX1_30/a_66_6# in_clkb DFFPOSX1_30/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5251 DFFPOSX1_30/a_76_6# DFFPOSX1_30/a_2_6# DFFPOSX1_30/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5252 gnd out_temp_addNum[0] DFFPOSX1_30/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5253 out_temp_addNum[0] DFFPOSX1_30/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5254 NOR2X1_13/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5255 NOR2X1_13/Y INVX2_59/Y NOR2X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5256 NOR2X1_13/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5257 gnd INVX2_59/Y NOR2X1_13/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5258 INVX2_46/Y INVX2_46/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5259 INVX2_46/Y INVX2_46/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5260 vdd BUFX2_0/A BUFX2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5261 BUFX2_1/Y BUFX2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5262 gnd BUFX2_0/A BUFX2_1/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M5263 BUFX2_1/Y BUFX2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5264 BUFX2_0/A in_clkb vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5265 BUFX2_0/A in_clkb gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5266 OAI21X1_37/a_9_54# INVX2_44/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5267 OAI21X1_44/C INVX2_46/Y OAI21X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5268 vdd con_readData OAI21X1_44/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5269 gnd INVX2_44/Y OAI21X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5270 OAI21X1_37/a_2_6# INVX2_46/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5271 OAI21X1_44/C con_readData OAI21X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5272 vdd BUFX2_0/A BUFX2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5273 BUFX2_0/Y BUFX2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5274 gnd BUFX2_0/A BUFX2_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M5275 BUFX2_0/Y BUFX2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5276 INVX2_43/Y BUFX2_0/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5277 INVX2_43/Y BUFX2_0/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5278 INVX2_41/Y BUFX2_0/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5279 INVX2_41/Y BUFX2_0/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5280 vdd INVX2_43/Y DFFPOSX1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5281 DFFPOSX1_29/a_17_74# OAI21X1_35/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5282 DFFPOSX1_29/a_22_6# INVX2_43/Y DFFPOSX1_29/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5283 DFFPOSX1_29/a_31_74# DFFPOSX1_29/a_2_6# DFFPOSX1_29/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5284 vdd DFFPOSX1_29/a_34_4# DFFPOSX1_29/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5285 DFFPOSX1_29/a_34_4# DFFPOSX1_29/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5286 DFFPOSX1_29/a_61_74# DFFPOSX1_29/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5287 DFFPOSX1_29/a_66_6# DFFPOSX1_29/a_2_6# DFFPOSX1_29/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5288 DFFPOSX1_29/a_76_84# INVX2_43/Y DFFPOSX1_29/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5289 vdd con_restart DFFPOSX1_29/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5290 gnd INVX2_43/Y DFFPOSX1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5291 con_restart DFFPOSX1_29/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5292 DFFPOSX1_29/a_17_6# OAI21X1_35/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5293 DFFPOSX1_29/a_22_6# DFFPOSX1_29/a_2_6# DFFPOSX1_29/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5294 DFFPOSX1_29/a_31_6# INVX2_43/Y DFFPOSX1_29/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5295 gnd DFFPOSX1_29/a_34_4# DFFPOSX1_29/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5296 DFFPOSX1_29/a_34_4# DFFPOSX1_29/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5297 DFFPOSX1_29/a_61_6# DFFPOSX1_29/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5298 DFFPOSX1_29/a_66_6# INVX2_43/Y DFFPOSX1_29/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5299 DFFPOSX1_29/a_76_6# DFFPOSX1_29/a_2_6# DFFPOSX1_29/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5300 gnd con_restart DFFPOSX1_29/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5301 con_restart DFFPOSX1_29/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5302 OAI21X1_35/a_9_54# BUFX2_2/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5303 OAI21X1_35/Y OAI21X1_35/B OAI21X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5304 vdd OAI21X1_52/C OAI21X1_35/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5305 gnd BUFX2_2/Y OAI21X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5306 OAI21X1_35/a_2_6# OAI21X1_35/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5307 OAI21X1_35/Y OAI21X1_52/C OAI21X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5308 vdd BUFX2_5/Y DFFPOSX1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5309 DFFPOSX1_27/a_17_74# NAND2X1_9/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5310 DFFPOSX1_27/a_22_6# BUFX2_5/Y DFFPOSX1_27/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5311 DFFPOSX1_27/a_31_74# DFFPOSX1_27/a_2_6# DFFPOSX1_27/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5312 vdd DFFPOSX1_27/a_34_4# DFFPOSX1_27/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5313 DFFPOSX1_27/a_34_4# DFFPOSX1_27/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5314 DFFPOSX1_27/a_61_74# DFFPOSX1_27/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5315 DFFPOSX1_27/a_66_6# DFFPOSX1_27/a_2_6# DFFPOSX1_27/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5316 DFFPOSX1_27/a_76_84# BUFX2_5/Y DFFPOSX1_27/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5317 vdd INVX2_51/A DFFPOSX1_27/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5318 gnd BUFX2_5/Y DFFPOSX1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5319 INVX2_51/A DFFPOSX1_27/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5320 DFFPOSX1_27/a_17_6# NAND2X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5321 DFFPOSX1_27/a_22_6# DFFPOSX1_27/a_2_6# DFFPOSX1_27/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5322 DFFPOSX1_27/a_31_6# BUFX2_5/Y DFFPOSX1_27/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5323 gnd DFFPOSX1_27/a_34_4# DFFPOSX1_27/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5324 DFFPOSX1_27/a_34_4# DFFPOSX1_27/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5325 DFFPOSX1_27/a_61_6# DFFPOSX1_27/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5326 DFFPOSX1_27/a_66_6# BUFX2_5/Y DFFPOSX1_27/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5327 DFFPOSX1_27/a_76_6# DFFPOSX1_27/a_2_6# DFFPOSX1_27/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5328 gnd INVX2_51/A DFFPOSX1_27/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5329 INVX2_51/A DFFPOSX1_27/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5330 INVX2_40/Y INVX2_40/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5331 INVX2_40/Y INVX2_40/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5332 vdd INVX2_43/Y DFFPOSX1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5333 DFFPOSX1_26/a_17_74# INVX2_51/A vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5334 DFFPOSX1_26/a_22_6# INVX2_43/Y DFFPOSX1_26/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5335 DFFPOSX1_26/a_31_74# DFFPOSX1_26/a_2_6# DFFPOSX1_26/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5336 vdd DFFPOSX1_26/a_34_4# DFFPOSX1_26/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5337 DFFPOSX1_26/a_34_4# DFFPOSX1_26/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5338 DFFPOSX1_26/a_61_74# DFFPOSX1_26/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5339 DFFPOSX1_26/a_66_6# DFFPOSX1_26/a_2_6# DFFPOSX1_26/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5340 DFFPOSX1_26/a_76_84# INVX2_43/Y DFFPOSX1_26/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5341 vdd out_state[0] DFFPOSX1_26/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5342 gnd INVX2_43/Y DFFPOSX1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5343 out_state[0] DFFPOSX1_26/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5344 DFFPOSX1_26/a_17_6# INVX2_51/A gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5345 DFFPOSX1_26/a_22_6# DFFPOSX1_26/a_2_6# DFFPOSX1_26/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5346 DFFPOSX1_26/a_31_6# INVX2_43/Y DFFPOSX1_26/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5347 gnd DFFPOSX1_26/a_34_4# DFFPOSX1_26/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5348 DFFPOSX1_26/a_34_4# DFFPOSX1_26/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5349 DFFPOSX1_26/a_61_6# DFFPOSX1_26/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5350 DFFPOSX1_26/a_66_6# INVX2_43/Y DFFPOSX1_26/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5351 DFFPOSX1_26/a_76_6# DFFPOSX1_26/a_2_6# DFFPOSX1_26/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5352 gnd out_state[0] DFFPOSX1_26/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5353 out_state[0] DFFPOSX1_26/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5354 vdd XOR2X1_50/A XOR2X1_50/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5355 XOR2X1_50/a_18_54# XOR2X1_50/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5356 XOR2X1_50/Y XOR2X1_50/A XOR2X1_50/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5357 XOR2X1_50/a_35_54# XOR2X1_50/a_2_6# XOR2X1_50/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5358 vdd XOR2X1_50/B XOR2X1_50/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5359 XOR2X1_50/a_13_43# XOR2X1_50/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5360 gnd XOR2X1_50/A XOR2X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5361 XOR2X1_50/a_18_6# XOR2X1_50/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5362 XOR2X1_50/Y XOR2X1_50/a_2_6# XOR2X1_50/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5363 XOR2X1_50/a_35_6# XOR2X1_50/A XOR2X1_50/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5364 gnd XOR2X1_50/B XOR2X1_50/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5365 XOR2X1_50/a_13_43# XOR2X1_50/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5366 NOR2X1_17/a_9_54# NOR2X1_17/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5367 NOR2X1_17/Y NOR2X1_17/B NOR2X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5368 NOR2X1_17/Y NOR2X1_17/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5369 gnd NOR2X1_17/B NOR2X1_17/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5370 vdd XNOR2X1_27/A XNOR2X1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5371 XNOR2X1_27/a_18_54# XNOR2X1_27/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5372 XNOR2X1_27/Y XNOR2X1_27/a_2_6# XNOR2X1_27/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5373 XNOR2X1_27/a_35_54# XNOR2X1_27/A XNOR2X1_27/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5374 vdd AND2X2_18/Y XNOR2X1_27/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5375 XNOR2X1_27/a_12_41# AND2X2_18/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5376 gnd XNOR2X1_27/A XNOR2X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5377 XNOR2X1_27/a_18_6# XNOR2X1_27/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5378 XNOR2X1_27/Y XNOR2X1_27/A XNOR2X1_27/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5379 XNOR2X1_27/a_35_6# XNOR2X1_27/a_2_6# XNOR2X1_27/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5380 gnd AND2X2_18/Y XNOR2X1_27/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5381 XNOR2X1_27/a_12_41# AND2X2_18/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5382 AND2X2_18/a_2_6# AND2X2_18/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5383 vdd AND2X2_18/B AND2X2_18/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5384 AND2X2_18/Y AND2X2_18/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5385 AND2X2_18/a_9_6# AND2X2_18/A AND2X2_18/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M5386 gnd AND2X2_18/B AND2X2_18/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5387 AND2X2_18/Y AND2X2_18/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5388 vdd INVX2_5/A XNOR2X1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5389 XNOR2X1_26/a_18_54# XNOR2X1_26/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5390 XOR2X1_48/B XNOR2X1_26/a_2_6# XNOR2X1_26/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5391 XNOR2X1_26/a_35_54# INVX2_5/A XOR2X1_48/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5392 vdd XOR2X1_52/Y XNOR2X1_26/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5393 XNOR2X1_26/a_12_41# XOR2X1_52/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5394 gnd INVX2_5/A XNOR2X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5395 XNOR2X1_26/a_18_6# XNOR2X1_26/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5396 XOR2X1_48/B INVX2_5/A XNOR2X1_26/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5397 XNOR2X1_26/a_35_6# XNOR2X1_26/a_2_6# XOR2X1_48/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5398 gnd XOR2X1_52/Y XNOR2X1_26/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5399 XNOR2X1_26/a_12_41# XOR2X1_52/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5400 NOR2X1_15/A AOI22X1_44/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5401 vdd NAND3X1_17/B NOR2X1_15/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5402 NOR2X1_15/A AND2X2_39/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5403 NAND3X1_17/a_9_6# AOI22X1_44/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5404 NAND3X1_17/a_14_6# NAND3X1_17/B NAND3X1_17/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5405 NOR2X1_15/A AND2X2_39/Y NAND3X1_17/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5406 OAI21X1_40/A NAND3X1_16/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5407 vdd NAND3X1_16/B OAI21X1_40/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5408 OAI21X1_40/A AND2X2_38/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5409 NAND3X1_16/a_9_6# NAND3X1_16/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5410 NAND3X1_16/a_14_6# NAND3X1_16/B NAND3X1_16/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5411 OAI21X1_40/A AND2X2_38/Y NAND3X1_16/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5412 INVX2_50/Y out_MuxData[13] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5413 INVX2_50/Y out_MuxData[13] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5414 vdd INVX2_5/A XOR2X1_46/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5415 XOR2X1_46/a_18_54# XOR2X1_46/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5416 XOR2X1_46/Y INVX2_5/A XOR2X1_46/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5417 XOR2X1_46/a_35_54# XOR2X1_46/a_2_6# XOR2X1_46/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5418 vdd XOR2X1_69/B XOR2X1_46/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5419 XOR2X1_46/a_13_43# XOR2X1_69/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5420 gnd INVX2_5/A XOR2X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5421 XOR2X1_46/a_18_6# XOR2X1_46/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5422 XOR2X1_46/Y XOR2X1_46/a_2_6# XOR2X1_46/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5423 XOR2X1_46/a_35_6# INVX2_5/A XOR2X1_46/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5424 gnd XOR2X1_69/B XOR2X1_46/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5425 XOR2X1_46/a_13_43# XOR2X1_69/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5426 vdd out_MuxData[9] AOI22X1_41/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5427 AOI22X1_41/a_2_54# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5428 AOI22X1_41/Y out_MuxData[13] AOI22X1_41/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5429 AOI22X1_41/a_2_54# XOR2X1_38/Y AOI22X1_41/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5430 AOI22X1_41/a_11_6# out_MuxData[9] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5431 AOI22X1_41/Y out_MuxData[7] AOI22X1_41/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5432 AOI22X1_41/a_28_6# out_MuxData[13] AOI22X1_41/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5433 gnd XOR2X1_38/Y AOI22X1_41/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5434 NOR2X1_15/a_9_54# NOR2X1_15/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5435 INVX2_44/A NOR2X1_15/B NOR2X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5436 INVX2_44/A NOR2X1_15/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5437 gnd NOR2X1_15/B INVX2_44/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5438 vdd XOR2X1_37/B AOI22X1_40/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5439 AOI22X1_40/a_2_54# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5440 NOR2X1_14/A out_MuxData[4] AOI22X1_40/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5441 AOI22X1_40/a_2_54# XOR2X1_36/B NOR2X1_14/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5442 AOI22X1_40/a_11_6# XOR2X1_37/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5443 NOR2X1_14/A out_MuxData[5] AOI22X1_40/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5444 AOI22X1_40/a_28_6# out_MuxData[4] NOR2X1_14/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5445 gnd XOR2X1_36/B AOI22X1_40/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5446 vdd NOR2X1_14/B XNOR2X1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5447 XNOR2X1_24/a_18_54# XNOR2X1_24/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5448 XNOR2X1_24/Y XNOR2X1_24/a_2_6# XNOR2X1_24/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5449 XNOR2X1_24/a_35_54# NOR2X1_14/B XNOR2X1_24/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5450 vdd NOR2X1_14/A XNOR2X1_24/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5451 XNOR2X1_24/a_12_41# NOR2X1_14/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5452 gnd NOR2X1_14/B XNOR2X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5453 XNOR2X1_24/a_18_6# XNOR2X1_24/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5454 XNOR2X1_24/Y NOR2X1_14/B XNOR2X1_24/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5455 XNOR2X1_24/a_35_6# XNOR2X1_24/a_2_6# XNOR2X1_24/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5456 gnd NOR2X1_14/A XNOR2X1_24/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5457 XNOR2X1_24/a_12_41# NOR2X1_14/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5458 INVX2_48/Y INVX2_48/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5459 INVX2_48/Y INVX2_48/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5460 vdd in_clkb DFFPOSX1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5461 DFFPOSX1_32/a_17_74# OAI22X1_1/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5462 DFFPOSX1_32/a_22_6# in_clkb DFFPOSX1_32/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5463 DFFPOSX1_32/a_31_74# DFFPOSX1_32/a_2_6# DFFPOSX1_32/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5464 vdd DFFPOSX1_32/a_34_4# DFFPOSX1_32/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5465 DFFPOSX1_32/a_34_4# DFFPOSX1_32/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5466 DFFPOSX1_32/a_61_74# DFFPOSX1_32/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5467 DFFPOSX1_32/a_66_6# DFFPOSX1_32/a_2_6# DFFPOSX1_32/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5468 DFFPOSX1_32/a_76_84# in_clkb DFFPOSX1_32/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5469 vdd INVX2_48/A DFFPOSX1_32/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5470 gnd in_clkb DFFPOSX1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5471 INVX2_48/A DFFPOSX1_32/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5472 DFFPOSX1_32/a_17_6# OAI22X1_1/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5473 DFFPOSX1_32/a_22_6# DFFPOSX1_32/a_2_6# DFFPOSX1_32/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5474 DFFPOSX1_32/a_31_6# in_clkb DFFPOSX1_32/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5475 gnd DFFPOSX1_32/a_34_4# DFFPOSX1_32/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5476 DFFPOSX1_32/a_34_4# DFFPOSX1_32/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5477 DFFPOSX1_32/a_61_6# DFFPOSX1_32/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5478 DFFPOSX1_32/a_66_6# in_clkb DFFPOSX1_32/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5479 DFFPOSX1_32/a_76_6# DFFPOSX1_32/a_2_6# DFFPOSX1_32/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5480 gnd INVX2_48/A DFFPOSX1_32/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5481 INVX2_48/A DFFPOSX1_32/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5482 OAI22X1_1/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5483 OAI22X1_1/Y INVX2_48/Y OAI22X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M5484 OAI22X1_1/a_28_54# INVX2_37/Y OAI22X1_1/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5485 vdd INVX2_62/Y OAI22X1_1/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5486 gnd BUFX2_3/Y OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M5487 OAI22X1_1/a_2_6# INVX2_48/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5488 OAI22X1_1/Y INVX2_37/Y OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5489 OAI22X1_1/a_2_6# INVX2_62/Y OAI22X1_1/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5490 OAI21X1_41/a_9_54# OAI21X1_40/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5491 OAI21X1_39/C NAND3X1_7/Y OAI21X1_41/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5492 vdd BUFX2_4/Y OAI21X1_39/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5493 gnd OAI21X1_40/A OAI21X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5494 OAI21X1_41/a_2_6# NAND3X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5495 OAI21X1_39/C BUFX2_4/Y OAI21X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5496 OAI21X1_40/a_9_54# OAI21X1_40/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5497 AOI22X1_38/A NAND3X1_7/Y OAI21X1_40/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5498 vdd INVX2_44/A AOI22X1_38/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5499 gnd OAI21X1_40/A OAI21X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5500 OAI21X1_40/a_2_6# NAND3X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5501 AOI22X1_38/A INVX2_44/A OAI21X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5502 OAI21X1_39/a_9_54# BUFX2_2/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5503 OAI21X1_39/Y INVX2_47/Y OAI21X1_39/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5504 vdd OAI21X1_39/C OAI21X1_39/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5505 gnd BUFX2_2/Y OAI21X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5506 OAI21X1_39/a_2_6# INVX2_47/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5507 OAI21X1_39/Y OAI21X1_39/C OAI21X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5508 INVX2_47/Y out_temp_addNum[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5509 INVX2_47/Y out_temp_addNum[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5510 OAI21X1_38/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5511 OAI21X1_38/Y INVX2_46/A OAI21X1_38/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5512 vdd OAI21X1_38/C OAI21X1_38/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5513 gnd con_restart OAI21X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5514 OAI21X1_38/a_2_6# INVX2_46/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5515 OAI21X1_38/Y OAI21X1_38/C OAI21X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5516 vdd AOI22X1_38/A AOI22X1_38/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5517 AOI22X1_38/a_2_54# INVX2_46/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5518 OAI22X1_3/C INVX2_44/A AOI22X1_38/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5519 AOI22X1_38/a_2_54# INVX2_46/A OAI22X1_3/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5520 AOI22X1_38/a_11_6# AOI22X1_38/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5521 OAI22X1_3/C INVX2_46/Y AOI22X1_38/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5522 AOI22X1_38/a_28_6# INVX2_44/A OAI22X1_3/C Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5523 gnd INVX2_46/A AOI22X1_38/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5524 INVX2_44/Y INVX2_44/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5525 INVX2_44/Y INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5526 INVX2_42/Y INVX2_42/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5527 INVX2_42/Y INVX2_42/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5528 OAI21X1_36/a_9_54# con_loseSig vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5529 INVX2_42/A INVX2_57/Y OAI21X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5530 vdd BUFX2_3/Y INVX2_42/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5531 gnd con_loseSig OAI21X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5532 OAI21X1_36/a_2_6# INVX2_57/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5533 INVX2_42/A BUFX2_3/Y OAI21X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5534 vdd BUFX2_9/Y DFFPOSX1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5535 DFFPOSX1_28/a_17_74# NAND2X1_11/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5536 DFFPOSX1_28/a_22_6# BUFX2_9/Y DFFPOSX1_28/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5537 DFFPOSX1_28/a_31_74# DFFPOSX1_28/a_2_6# DFFPOSX1_28/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5538 vdd DFFPOSX1_28/a_34_4# DFFPOSX1_28/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5539 DFFPOSX1_28/a_34_4# DFFPOSX1_28/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5540 DFFPOSX1_28/a_61_74# DFFPOSX1_28/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5541 DFFPOSX1_28/a_66_6# DFFPOSX1_28/a_2_6# DFFPOSX1_28/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5542 DFFPOSX1_28/a_76_84# BUFX2_9/Y DFFPOSX1_28/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5543 vdd INVX2_40/A DFFPOSX1_28/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5544 gnd BUFX2_9/Y DFFPOSX1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5545 INVX2_40/A DFFPOSX1_28/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5546 DFFPOSX1_28/a_17_6# NAND2X1_11/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5547 DFFPOSX1_28/a_22_6# DFFPOSX1_28/a_2_6# DFFPOSX1_28/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5548 DFFPOSX1_28/a_31_6# BUFX2_9/Y DFFPOSX1_28/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5549 gnd DFFPOSX1_28/a_34_4# DFFPOSX1_28/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5550 DFFPOSX1_28/a_34_4# DFFPOSX1_28/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5551 DFFPOSX1_28/a_61_6# DFFPOSX1_28/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5552 DFFPOSX1_28/a_66_6# BUFX2_9/Y DFFPOSX1_28/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5553 DFFPOSX1_28/a_76_6# DFFPOSX1_28/a_2_6# DFFPOSX1_28/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5554 gnd INVX2_40/A DFFPOSX1_28/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5555 INVX2_40/A DFFPOSX1_28/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5556 OAI21X1_35/B INVX2_11/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5557 vdd INVX2_53/A OAI21X1_35/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5558 NAND2X1_15/a_9_6# INVX2_11/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5559 OAI21X1_35/B INVX2_53/A NAND2X1_15/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5560 vdd BUFX2_5/Y DFFPOSX1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5561 DFFPOSX1_25/a_17_74# NAND3X1_12/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5562 DFFPOSX1_25/a_22_6# BUFX2_5/Y DFFPOSX1_25/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5563 DFFPOSX1_25/a_31_74# DFFPOSX1_25/a_2_6# DFFPOSX1_25/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5564 vdd DFFPOSX1_25/a_34_4# DFFPOSX1_25/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5565 DFFPOSX1_25/a_34_4# DFFPOSX1_25/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5566 DFFPOSX1_25/a_61_74# DFFPOSX1_25/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5567 DFFPOSX1_25/a_66_6# DFFPOSX1_25/a_2_6# DFFPOSX1_25/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5568 DFFPOSX1_25/a_76_84# BUFX2_5/Y DFFPOSX1_25/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5569 vdd INVX2_52/A DFFPOSX1_25/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5570 gnd BUFX2_5/Y DFFPOSX1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5571 INVX2_52/A DFFPOSX1_25/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5572 DFFPOSX1_25/a_17_6# NAND3X1_12/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5573 DFFPOSX1_25/a_22_6# DFFPOSX1_25/a_2_6# DFFPOSX1_25/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5574 DFFPOSX1_25/a_31_6# BUFX2_5/Y DFFPOSX1_25/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5575 gnd DFFPOSX1_25/a_34_4# DFFPOSX1_25/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5576 DFFPOSX1_25/a_34_4# DFFPOSX1_25/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5577 DFFPOSX1_25/a_61_6# DFFPOSX1_25/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5578 DFFPOSX1_25/a_66_6# BUFX2_5/Y DFFPOSX1_25/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5579 DFFPOSX1_25/a_76_6# DFFPOSX1_25/a_2_6# DFFPOSX1_25/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5580 gnd INVX2_52/A DFFPOSX1_25/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5581 INVX2_52/A DFFPOSX1_25/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5582 vdd INVX2_43/Y DFFPOSX1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5583 DFFPOSX1_24/a_17_74# INVX2_52/A vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5584 DFFPOSX1_24/a_22_6# INVX2_43/Y DFFPOSX1_24/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5585 DFFPOSX1_24/a_31_74# DFFPOSX1_24/a_2_6# DFFPOSX1_24/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5586 vdd DFFPOSX1_24/a_34_4# DFFPOSX1_24/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5587 DFFPOSX1_24/a_34_4# DFFPOSX1_24/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5588 DFFPOSX1_24/a_61_74# DFFPOSX1_24/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5589 DFFPOSX1_24/a_66_6# DFFPOSX1_24/a_2_6# DFFPOSX1_24/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5590 DFFPOSX1_24/a_76_84# INVX2_43/Y DFFPOSX1_24/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5591 vdd out_state[1] DFFPOSX1_24/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5592 gnd INVX2_43/Y DFFPOSX1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5593 out_state[1] DFFPOSX1_24/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5594 DFFPOSX1_24/a_17_6# INVX2_52/A gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5595 DFFPOSX1_24/a_22_6# DFFPOSX1_24/a_2_6# DFFPOSX1_24/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5596 DFFPOSX1_24/a_31_6# INVX2_43/Y DFFPOSX1_24/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5597 gnd DFFPOSX1_24/a_34_4# DFFPOSX1_24/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5598 DFFPOSX1_24/a_34_4# DFFPOSX1_24/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5599 DFFPOSX1_24/a_61_6# DFFPOSX1_24/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5600 DFFPOSX1_24/a_66_6# INVX2_43/Y DFFPOSX1_24/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5601 DFFPOSX1_24/a_76_6# DFFPOSX1_24/a_2_6# DFFPOSX1_24/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5602 gnd out_state[1] DFFPOSX1_24/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5603 out_state[1] DFFPOSX1_24/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5604 OAI21X1_34/a_9_54# AOI22X1_36/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5605 XOR2X1_50/A OAI21X1_33/B OAI21X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5606 vdd NAND3X1_15/Y XOR2X1_50/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5607 gnd AOI22X1_36/Y OAI21X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5608 OAI21X1_34/a_2_6# OAI21X1_33/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5609 XOR2X1_50/A NAND3X1_15/Y OAI21X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5610 NAND3X1_15/B AOI22X1_36/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5611 vdd OAI21X1_33/B NAND3X1_15/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5612 NAND2X1_14/a_9_6# AOI22X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5613 NAND3X1_15/B OAI21X1_33/B NAND2X1_14/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5614 OAI21X1_33/a_9_54# AOI22X1_36/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5615 XNOR2X1_27/A OAI21X1_33/B OAI21X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5616 vdd NAND3X1_15/B XNOR2X1_27/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5617 gnd AOI22X1_36/Y OAI21X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5618 OAI21X1_33/a_2_6# OAI21X1_33/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5619 XNOR2X1_27/A NAND3X1_15/B OAI21X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5620 NAND3X1_15/Y AND2X2_18/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5621 vdd NAND3X1_15/B NAND3X1_15/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5622 NAND3X1_15/Y AND2X2_18/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5623 NAND3X1_15/a_9_6# AND2X2_18/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5624 NAND3X1_15/a_14_6# NAND3X1_15/B NAND3X1_15/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5625 NAND3X1_15/Y AND2X2_18/B NAND3X1_15/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5626 vdd AND2X2_18/B XOR2X1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5627 XOR2X1_44/a_18_54# XOR2X1_44/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5628 XOR2X1_44/Y AND2X2_18/B XOR2X1_44/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5629 XOR2X1_44/a_35_54# XOR2X1_44/a_2_6# XOR2X1_44/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5630 vdd AND2X2_18/A XOR2X1_44/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5631 XOR2X1_44/a_13_43# AND2X2_18/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5632 gnd AND2X2_18/B XOR2X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5633 XOR2X1_44/a_18_6# XOR2X1_44/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5634 XOR2X1_44/Y XOR2X1_44/a_2_6# XOR2X1_44/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5635 XOR2X1_44/a_35_6# AND2X2_18/B XOR2X1_44/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5636 gnd AND2X2_18/A XOR2X1_44/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5637 XOR2X1_44/a_13_43# AND2X2_18/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5638 vdd out_MuxData[3] AOI22X1_36/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5639 AOI22X1_36/a_2_54# out_MuxData[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5640 AOI22X1_36/Y out_MuxData[7] AOI22X1_36/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5641 AOI22X1_36/a_2_54# XOR2X1_47/Y AOI22X1_36/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5642 AOI22X1_36/a_11_6# out_MuxData[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5643 AOI22X1_36/Y out_MuxData[13] AOI22X1_36/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5644 AOI22X1_36/a_28_6# out_MuxData[7] AOI22X1_36/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5645 gnd XOR2X1_47/Y AOI22X1_36/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5646 AND2X2_17/a_2_6# AND2X2_17/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5647 vdd AND2X2_17/B AND2X2_17/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5648 AND2X2_17/Y AND2X2_17/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5649 AND2X2_17/a_9_6# AND2X2_17/A AND2X2_17/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M5650 gnd AND2X2_17/B AND2X2_17/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5651 AND2X2_17/Y AND2X2_17/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5652 vdd INVX2_17/Y XNOR2X1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5653 XNOR2X1_20/a_18_54# XNOR2X1_20/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5654 AND2X2_18/B XNOR2X1_20/a_2_6# XNOR2X1_20/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5655 XNOR2X1_20/a_35_54# INVX2_17/Y AND2X2_18/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5656 vdd XOR2X1_47/Y XNOR2X1_20/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5657 XNOR2X1_20/a_12_41# XOR2X1_47/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5658 gnd INVX2_17/Y XNOR2X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5659 XNOR2X1_20/a_18_6# XNOR2X1_20/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5660 AND2X2_18/B INVX2_17/Y XNOR2X1_20/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5661 XNOR2X1_20/a_35_6# XNOR2X1_20/a_2_6# AND2X2_18/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5662 gnd XOR2X1_47/Y XNOR2X1_20/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5663 XNOR2X1_20/a_12_41# XOR2X1_47/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5664 vdd AOI22X1_35/A AOI22X1_35/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5665 AOI22X1_35/a_2_54# INVX2_71/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5666 AND2X2_17/B INVX2_59/Y AOI22X1_35/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5667 AOI22X1_35/a_2_54# XNOR2X1_27/Y AND2X2_17/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5668 AOI22X1_35/a_11_6# AOI22X1_35/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5669 AND2X2_17/B INVX2_71/Y AOI22X1_35/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5670 AOI22X1_35/a_28_6# INVX2_59/Y AND2X2_17/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5671 gnd XNOR2X1_27/Y AOI22X1_35/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5672 vdd INVX2_59/Y AOI22X1_34/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5673 AOI22X1_34/a_2_54# XOR2X1_44/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5674 NAND3X1_16/A XOR2X1_40/Y AOI22X1_34/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5675 AOI22X1_34/a_2_54# INVX2_71/Y NAND3X1_16/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5676 AOI22X1_34/a_11_6# INVX2_59/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5677 NAND3X1_16/A XOR2X1_44/Y AOI22X1_34/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5678 AOI22X1_34/a_28_6# XOR2X1_40/Y NAND3X1_16/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5679 gnd INVX2_71/Y AOI22X1_34/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5680 INVX2_5/A INVX2_39/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5681 INVX2_5/A INVX2_39/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5682 vdd INVX2_17/Y XOR2X1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5683 XOR2X1_38/a_18_54# XOR2X1_38/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5684 XOR2X1_38/Y INVX2_17/Y XOR2X1_38/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5685 XOR2X1_38/a_35_54# XOR2X1_38/a_2_6# XOR2X1_38/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5686 vdd XOR2X1_69/B XOR2X1_38/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5687 XOR2X1_38/a_13_43# XOR2X1_69/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5688 gnd INVX2_17/Y XOR2X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5689 XOR2X1_38/a_18_6# XOR2X1_38/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5690 XOR2X1_38/Y XOR2X1_38/a_2_6# XOR2X1_38/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5691 XOR2X1_38/a_35_6# INVX2_17/Y XOR2X1_38/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5692 gnd XOR2X1_69/B XOR2X1_38/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5693 XOR2X1_38/a_13_43# XOR2X1_69/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5694 vdd INVX2_50/Y XNOR2X1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5695 XNOR2X1_18/a_18_54# XNOR2X1_18/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5696 XOR2X1_33/B XNOR2X1_18/a_2_6# XNOR2X1_18/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5697 XNOR2X1_18/a_35_54# INVX2_50/Y XOR2X1_33/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5698 vdd XOR2X1_38/Y XNOR2X1_18/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5699 XNOR2X1_18/a_12_41# XOR2X1_38/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5700 gnd INVX2_50/Y XNOR2X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5701 XNOR2X1_18/a_18_6# XNOR2X1_18/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5702 XOR2X1_33/B INVX2_50/Y XNOR2X1_18/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5703 XNOR2X1_18/a_35_6# XNOR2X1_18/a_2_6# XOR2X1_33/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5704 gnd XOR2X1_38/Y XNOR2X1_18/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5705 XNOR2X1_18/a_12_41# XOR2X1_38/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5706 NOR2X1_15/B NAND3X1_14/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5707 vdd AOI22X1_30/Y NOR2X1_15/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5708 NOR2X1_15/B AND2X2_20/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5709 NAND3X1_14/a_9_6# NAND3X1_14/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5710 NAND3X1_14/a_14_6# AOI22X1_30/Y NAND3X1_14/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5711 NOR2X1_15/B AND2X2_20/Y NAND3X1_14/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5712 vdd out_MuxData[5] XOR2X1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5713 XOR2X1_37/a_18_54# XOR2X1_37/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5714 XOR2X1_36/B out_MuxData[5] XOR2X1_37/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5715 XOR2X1_37/a_35_54# XOR2X1_37/a_2_6# XOR2X1_36/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5716 vdd XOR2X1_37/B XOR2X1_37/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5717 XOR2X1_37/a_13_43# XOR2X1_37/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5718 gnd out_MuxData[5] XOR2X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5719 XOR2X1_37/a_18_6# XOR2X1_37/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5720 XOR2X1_36/B XOR2X1_37/a_2_6# XOR2X1_37/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5721 XOR2X1_37/a_35_6# out_MuxData[5] XOR2X1_36/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5722 gnd XOR2X1_37/B XOR2X1_37/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5723 XOR2X1_37/a_13_43# XOR2X1_37/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5724 vdd out_MuxData[4] XOR2X1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5725 XOR2X1_36/a_18_54# XOR2X1_36/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5726 XOR2X1_33/A out_MuxData[4] XOR2X1_36/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5727 XOR2X1_36/a_35_54# XOR2X1_36/a_2_6# XOR2X1_33/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5728 vdd XOR2X1_36/B XOR2X1_36/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5729 XOR2X1_36/a_13_43# XOR2X1_36/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5730 gnd out_MuxData[4] XOR2X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5731 XOR2X1_36/a_18_6# XOR2X1_36/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5732 XOR2X1_33/A XOR2X1_36/a_2_6# XOR2X1_36/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5733 XOR2X1_36/a_35_6# out_MuxData[4] XOR2X1_33/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5734 gnd XOR2X1_36/B XOR2X1_36/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5735 XOR2X1_36/a_13_43# XOR2X1_36/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5736 OAI21X1_32/a_9_54# AOI22X1_41/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5737 XOR2X1_34/A XNOR2X1_24/Y OAI21X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5738 vdd OAI21X1_32/C XOR2X1_34/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5739 gnd AOI22X1_41/Y OAI21X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5740 OAI21X1_32/a_2_6# XNOR2X1_24/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5741 XOR2X1_34/A OAI21X1_32/C OAI21X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5742 vdd XOR2X1_34/A XOR2X1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5743 XOR2X1_34/a_18_54# XOR2X1_34/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5744 XOR2X1_34/Y XOR2X1_34/A XOR2X1_34/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5745 XOR2X1_34/a_35_54# XOR2X1_34/a_2_6# XOR2X1_34/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5746 vdd NOR2X1_14/Y XOR2X1_34/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5747 XOR2X1_34/a_13_43# NOR2X1_14/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5748 gnd XOR2X1_34/A XOR2X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5749 XOR2X1_34/a_18_6# XOR2X1_34/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5750 XOR2X1_34/Y XOR2X1_34/a_2_6# XOR2X1_34/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5751 XOR2X1_34/a_35_6# XOR2X1_34/A XOR2X1_34/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5752 gnd NOR2X1_14/Y XOR2X1_34/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5753 XOR2X1_34/a_13_43# NOR2X1_14/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5754 vdd INVX2_104/Y AOI22X1_30/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5755 AOI22X1_30/a_2_54# XOR2X1_34/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5756 AOI22X1_30/Y XOR2X1_0/Y AOI22X1_30/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5757 AOI22X1_30/a_2_54# NOR2X1_41/B AOI22X1_30/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5758 AOI22X1_30/a_11_6# INVX2_104/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5759 AOI22X1_30/Y XOR2X1_34/Y AOI22X1_30/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5760 AOI22X1_30/a_28_6# XOR2X1_0/Y AOI22X1_30/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5761 gnd NOR2X1_41/B AOI22X1_30/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5762 INVX2_38/Y out_MemBData[3] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5763 INVX2_38/Y out_MemBData[3] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5764 OAI21X1_31/a_9_54# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5765 OAI21X1_31/Y OR2X2_0/Y OAI21X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5766 vdd OAI21X1_31/C OAI21X1_31/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5767 gnd INVX2_26/A OAI21X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5768 OAI21X1_31/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5769 OAI21X1_31/Y OAI21X1_31/C OAI21X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5770 INVX2_37/Y out_MemBData[1] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5771 INVX2_37/Y out_MemBData[1] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5772 vdd BUFX2_11/Y DFFPOSX1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5773 DFFPOSX1_22/a_17_74# OAI21X1_30/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5774 DFFPOSX1_22/a_22_6# BUFX2_11/Y DFFPOSX1_22/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5775 DFFPOSX1_22/a_31_74# DFFPOSX1_22/a_2_6# DFFPOSX1_22/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5776 vdd DFFPOSX1_22/a_34_4# DFFPOSX1_22/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5777 DFFPOSX1_22/a_34_4# DFFPOSX1_22/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5778 DFFPOSX1_22/a_61_74# DFFPOSX1_22/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5779 DFFPOSX1_22/a_66_6# DFFPOSX1_22/a_2_6# DFFPOSX1_22/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5780 DFFPOSX1_22/a_76_84# BUFX2_11/Y DFFPOSX1_22/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5781 vdd out_MemBData[1] DFFPOSX1_22/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5782 gnd BUFX2_11/Y DFFPOSX1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5783 out_MemBData[1] DFFPOSX1_22/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5784 DFFPOSX1_22/a_17_6# OAI21X1_30/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5785 DFFPOSX1_22/a_22_6# DFFPOSX1_22/a_2_6# DFFPOSX1_22/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5786 DFFPOSX1_22/a_31_6# BUFX2_11/Y DFFPOSX1_22/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5787 gnd DFFPOSX1_22/a_34_4# DFFPOSX1_22/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5788 DFFPOSX1_22/a_34_4# DFFPOSX1_22/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5789 DFFPOSX1_22/a_61_6# DFFPOSX1_22/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5790 DFFPOSX1_22/a_66_6# BUFX2_11/Y DFFPOSX1_22/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5791 DFFPOSX1_22/a_76_6# DFFPOSX1_22/a_2_6# DFFPOSX1_22/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5792 gnd out_MemBData[1] DFFPOSX1_22/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5793 out_MemBData[1] DFFPOSX1_22/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5794 vdd in_clkb DFFPOSX1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5795 DFFPOSX1_21/a_17_74# OAI21X1_38/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5796 DFFPOSX1_21/a_22_6# in_clkb DFFPOSX1_21/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5797 DFFPOSX1_21/a_31_74# DFFPOSX1_21/a_2_6# DFFPOSX1_21/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5798 vdd DFFPOSX1_21/a_34_4# DFFPOSX1_21/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5799 DFFPOSX1_21/a_34_4# DFFPOSX1_21/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5800 DFFPOSX1_21/a_61_74# DFFPOSX1_21/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5801 DFFPOSX1_21/a_66_6# DFFPOSX1_21/a_2_6# DFFPOSX1_21/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5802 DFFPOSX1_21/a_76_84# in_clkb DFFPOSX1_21/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5803 vdd out_temp_addNum[1] DFFPOSX1_21/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5804 gnd in_clkb DFFPOSX1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5805 out_temp_addNum[1] DFFPOSX1_21/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5806 DFFPOSX1_21/a_17_6# OAI21X1_38/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5807 DFFPOSX1_21/a_22_6# DFFPOSX1_21/a_2_6# DFFPOSX1_21/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5808 DFFPOSX1_21/a_31_6# in_clkb DFFPOSX1_21/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5809 gnd DFFPOSX1_21/a_34_4# DFFPOSX1_21/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5810 DFFPOSX1_21/a_34_4# DFFPOSX1_21/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5811 DFFPOSX1_21/a_61_6# DFFPOSX1_21/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5812 DFFPOSX1_21/a_66_6# in_clkb DFFPOSX1_21/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5813 DFFPOSX1_21/a_76_6# DFFPOSX1_21/a_2_6# DFFPOSX1_21/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5814 gnd out_temp_addNum[1] DFFPOSX1_21/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5815 out_temp_addNum[1] DFFPOSX1_21/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5816 OAI21X1_38/C out_temp_addNum[1] vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5817 vdd con_restart OAI21X1_38/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5818 NAND2X1_12/a_9_6# out_temp_addNum[1] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5819 OAI21X1_38/C con_restart NAND2X1_12/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5820 vdd INVX2_41/Y DFFPOSX1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5821 DFFPOSX1_20/a_17_74# INVX2_42/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5822 DFFPOSX1_20/a_22_6# INVX2_41/Y DFFPOSX1_20/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5823 DFFPOSX1_20/a_31_74# DFFPOSX1_20/a_2_6# DFFPOSX1_20/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5824 vdd DFFPOSX1_20/a_34_4# DFFPOSX1_20/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5825 DFFPOSX1_20/a_34_4# DFFPOSX1_20/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5826 DFFPOSX1_20/a_61_74# DFFPOSX1_20/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5827 DFFPOSX1_20/a_66_6# DFFPOSX1_20/a_2_6# DFFPOSX1_20/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5828 DFFPOSX1_20/a_76_84# INVX2_41/Y DFFPOSX1_20/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5829 vdd con_loseSig DFFPOSX1_20/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5830 gnd INVX2_41/Y DFFPOSX1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5831 con_loseSig DFFPOSX1_20/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5832 DFFPOSX1_20/a_17_6# INVX2_42/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5833 DFFPOSX1_20/a_22_6# DFFPOSX1_20/a_2_6# DFFPOSX1_20/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5834 DFFPOSX1_20/a_31_6# INVX2_41/Y DFFPOSX1_20/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5835 gnd DFFPOSX1_20/a_34_4# DFFPOSX1_20/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5836 DFFPOSX1_20/a_34_4# DFFPOSX1_20/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5837 DFFPOSX1_20/a_61_6# DFFPOSX1_20/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5838 DFFPOSX1_20/a_66_6# INVX2_41/Y DFFPOSX1_20/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5839 DFFPOSX1_20/a_76_6# DFFPOSX1_20/a_2_6# DFFPOSX1_20/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5840 gnd con_loseSig DFFPOSX1_20/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5841 con_loseSig DFFPOSX1_20/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5842 vdd INVX2_41/Y DFFPOSX1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5843 DFFPOSX1_19/a_17_74# INVX2_40/A vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5844 DFFPOSX1_19/a_22_6# INVX2_41/Y DFFPOSX1_19/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5845 DFFPOSX1_19/a_31_74# DFFPOSX1_19/a_2_6# DFFPOSX1_19/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M5846 vdd DFFPOSX1_19/a_34_4# DFFPOSX1_19/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5847 DFFPOSX1_19/a_34_4# DFFPOSX1_19/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5848 DFFPOSX1_19/a_61_74# DFFPOSX1_19/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5849 DFFPOSX1_19/a_66_6# DFFPOSX1_19/a_2_6# DFFPOSX1_19/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M5850 DFFPOSX1_19/a_76_84# INVX2_41/Y DFFPOSX1_19/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5851 vdd out_state[2] DFFPOSX1_19/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5852 gnd INVX2_41/Y DFFPOSX1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5853 out_state[2] DFFPOSX1_19/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5854 DFFPOSX1_19/a_17_6# INVX2_40/A gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5855 DFFPOSX1_19/a_22_6# DFFPOSX1_19/a_2_6# DFFPOSX1_19/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5856 DFFPOSX1_19/a_31_6# INVX2_41/Y DFFPOSX1_19/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5857 gnd DFFPOSX1_19/a_34_4# DFFPOSX1_19/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5858 DFFPOSX1_19/a_34_4# DFFPOSX1_19/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M5859 DFFPOSX1_19/a_61_6# DFFPOSX1_19/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5860 DFFPOSX1_19/a_66_6# INVX2_41/Y DFFPOSX1_19/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M5861 DFFPOSX1_19/a_76_6# DFFPOSX1_19/a_2_6# DFFPOSX1_19/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M5862 gnd out_state[2] DFFPOSX1_19/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5863 out_state[2] DFFPOSX1_19/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5864 NAND2X1_11/Y AOI21X1_5/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M5865 vdd AOI21X1_2/Y NAND2X1_11/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5866 NAND2X1_11/a_9_6# AOI21X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5867 NAND2X1_11/Y AOI21X1_2/Y NAND2X1_11/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5868 INVX2_35/Y INVX2_35/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5869 INVX2_35/Y INVX2_35/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5870 vdd NOR2X1_10/B AOI21X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M5871 AOI21X1_5/a_2_54# INVX2_34/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5872 AOI21X1_5/Y INVX2_35/A AOI21X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5873 AOI21X1_5/a_12_6# NOR2X1_10/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5874 AOI21X1_5/Y INVX2_34/Y AOI21X1_5/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M5875 gnd INVX2_35/A AOI21X1_5/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5876 INVX2_34/Y out_state[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5877 INVX2_34/Y out_state[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5878 NAND3X1_12/Y OAI21X1_27/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M5879 vdd NAND3X1_6/Y NAND3X1_12/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5880 NAND3X1_12/Y INVX2_35/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5881 NAND3X1_12/a_9_6# OAI21X1_27/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5882 NAND3X1_12/a_14_6# NAND3X1_6/Y NAND3X1_12/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M5883 NAND3X1_12/Y INVX2_35/Y NAND3X1_12/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M5884 OAI21X1_27/a_9_54# out_state[2] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5885 OAI21X1_27/Y INVX2_70/Y OAI21X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M5886 vdd out_state[1] OAI21X1_27/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5887 gnd out_state[2] OAI21X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M5888 OAI21X1_27/a_2_6# INVX2_70/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5889 OAI21X1_27/Y out_state[1] OAI21X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5890 NOR2X1_11/a_9_54# INVX2_32/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5891 NOR2X1_10/B INVX2_70/Y NOR2X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5892 NOR2X1_10/B INVX2_32/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5893 gnd INVX2_70/Y NOR2X1_10/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5894 NOR2X1_10/a_9_54# out_state[2] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5895 AOI21X1_4/A NOR2X1_10/B NOR2X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5896 AOI21X1_4/A out_state[2] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5897 gnd NOR2X1_10/B AOI21X1_4/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5898 vdd AOI21X1_4/A AOI21X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M5899 AOI21X1_4/a_2_54# out_state[0] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5900 AOI21X1_4/Y AOI21X1_4/C AOI21X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5901 AOI21X1_4/a_12_6# AOI21X1_4/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5902 AOI21X1_4/Y out_state[0] AOI21X1_4/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M5903 gnd AOI21X1_4/C AOI21X1_4/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5904 NOR2X1_12/a_9_54# NOR2X1_12/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5905 XOR2X1_50/B NOR2X1_12/B NOR2X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5906 XOR2X1_50/B NOR2X1_12/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M5907 gnd NOR2X1_12/B XOR2X1_50/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5908 vdd NOR2X1_12/B XNOR2X1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5909 XNOR2X1_23/a_18_54# XNOR2X1_23/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5910 OAI21X1_33/B XNOR2X1_23/a_2_6# XNOR2X1_23/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5911 XNOR2X1_23/a_35_54# NOR2X1_12/B OAI21X1_33/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5912 vdd NOR2X1_12/A XNOR2X1_23/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5913 XNOR2X1_23/a_12_41# NOR2X1_12/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5914 gnd NOR2X1_12/B XNOR2X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5915 XNOR2X1_23/a_18_6# XNOR2X1_23/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5916 OAI21X1_33/B NOR2X1_12/B XNOR2X1_23/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5917 XNOR2X1_23/a_35_6# XNOR2X1_23/a_2_6# OAI21X1_33/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5918 gnd NOR2X1_12/A XNOR2X1_23/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5919 XNOR2X1_23/a_12_41# NOR2X1_12/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5920 vdd out_MuxData[6] AOI22X1_37/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5921 AOI22X1_37/a_2_54# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5922 NOR2X1_12/B out_MuxData[1] AOI22X1_37/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5923 AOI22X1_37/a_2_54# XOR2X1_32/Y NOR2X1_12/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5924 AOI22X1_37/a_11_6# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5925 NOR2X1_12/B out_MuxData[5] AOI22X1_37/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5926 AOI22X1_37/a_28_6# out_MuxData[1] NOR2X1_12/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5927 gnd XOR2X1_32/Y AOI22X1_37/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5928 vdd XNOR2X1_22/A XNOR2X1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5929 XNOR2X1_22/a_18_54# XNOR2X1_22/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5930 XOR2X1_42/A XNOR2X1_22/a_2_6# XNOR2X1_22/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5931 XNOR2X1_22/a_35_54# XNOR2X1_22/A XOR2X1_42/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5932 vdd out_MuxData[1] XNOR2X1_22/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5933 XNOR2X1_22/a_12_41# out_MuxData[1] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5934 gnd XNOR2X1_22/A XNOR2X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5935 XNOR2X1_22/a_18_6# XNOR2X1_22/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5936 XOR2X1_42/A XNOR2X1_22/A XNOR2X1_22/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5937 XNOR2X1_22/a_35_6# XNOR2X1_22/a_2_6# XOR2X1_42/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5938 gnd out_MuxData[1] XNOR2X1_22/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5939 XNOR2X1_22/a_12_41# out_MuxData[1] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5940 vdd INVX2_28/Y XNOR2X1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5941 XNOR2X1_21/a_18_54# XNOR2X1_21/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5942 AND2X2_18/A XNOR2X1_21/a_2_6# XNOR2X1_21/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5943 XNOR2X1_21/a_35_54# INVX2_28/Y AND2X2_18/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5944 vdd XOR2X1_43/Y XNOR2X1_21/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5945 XNOR2X1_21/a_12_41# XOR2X1_43/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5946 gnd INVX2_28/Y XNOR2X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5947 XNOR2X1_21/a_18_6# XNOR2X1_21/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5948 AND2X2_18/A INVX2_28/Y XNOR2X1_21/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5949 XNOR2X1_21/a_35_6# XNOR2X1_21/a_2_6# AND2X2_18/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5950 gnd XOR2X1_43/Y XNOR2X1_21/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5951 XNOR2X1_21/a_12_41# XOR2X1_43/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5952 vdd INVX2_39/A XOR2X1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5953 XOR2X1_43/a_18_54# XOR2X1_43/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5954 XOR2X1_43/Y INVX2_39/A XOR2X1_43/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5955 XOR2X1_43/a_35_54# XOR2X1_43/a_2_6# XOR2X1_43/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5956 vdd XOR2X1_43/B XOR2X1_43/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5957 XOR2X1_43/a_13_43# XOR2X1_43/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5958 gnd INVX2_39/A XOR2X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5959 XOR2X1_43/a_18_6# XOR2X1_43/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5960 XOR2X1_43/Y XOR2X1_43/a_2_6# XOR2X1_43/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5961 XOR2X1_43/a_35_6# INVX2_39/A XOR2X1_43/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5962 gnd XOR2X1_43/B XOR2X1_43/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5963 XOR2X1_43/a_13_43# XOR2X1_43/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5964 vdd XOR2X1_42/A AOI22X1_33/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M5965 AOI22X1_33/a_2_54# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5966 NOR2X1_9/B out_MuxData[3] AOI22X1_33/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M5967 AOI22X1_33/a_2_54# XOR2X1_41/A NOR2X1_9/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5968 AOI22X1_33/a_11_6# XOR2X1_42/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5969 NOR2X1_9/B out_MuxData[7] AOI22X1_33/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5970 AOI22X1_33/a_28_6# out_MuxData[3] NOR2X1_9/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5971 gnd XOR2X1_41/A AOI22X1_33/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5972 vdd XOR2X1_42/A XOR2X1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5973 XOR2X1_42/a_18_54# XOR2X1_42/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5974 XOR2X1_41/A XOR2X1_42/A XOR2X1_42/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5975 XOR2X1_42/a_35_54# XOR2X1_42/a_2_6# XOR2X1_41/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5976 vdd out_MuxData[7] XOR2X1_42/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5977 XOR2X1_42/a_13_43# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5978 gnd XOR2X1_42/A XOR2X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5979 XOR2X1_42/a_18_6# XOR2X1_42/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5980 XOR2X1_41/A XOR2X1_42/a_2_6# XOR2X1_42/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5981 XOR2X1_42/a_35_6# XOR2X1_42/A XOR2X1_41/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5982 gnd out_MuxData[7] XOR2X1_42/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5983 XOR2X1_42/a_13_43# out_MuxData[7] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5984 vdd XOR2X1_41/A XOR2X1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5985 XOR2X1_41/a_18_54# XOR2X1_41/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5986 XOR2X1_40/A XOR2X1_41/A XOR2X1_41/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5987 XOR2X1_41/a_35_54# XOR2X1_41/a_2_6# XOR2X1_40/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5988 vdd INVX2_86/A XOR2X1_41/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5989 XOR2X1_41/a_13_43# INVX2_86/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M5990 gnd XOR2X1_41/A XOR2X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M5991 XOR2X1_41/a_18_6# XOR2X1_41/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5992 XOR2X1_40/A XOR2X1_41/a_2_6# XOR2X1_41/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M5993 XOR2X1_41/a_35_6# XOR2X1_41/A XOR2X1_40/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M5994 gnd INVX2_86/A XOR2X1_41/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5995 XOR2X1_41/a_13_43# INVX2_86/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M5996 vdd XNOR2X1_19/A XNOR2X1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M5997 XNOR2X1_19/a_18_54# XNOR2X1_19/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M5998 AOI22X1_35/A XNOR2X1_19/a_2_6# XNOR2X1_19/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M5999 XNOR2X1_19/a_35_54# XNOR2X1_19/A AOI22X1_35/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6000 vdd AND2X2_16/Y XNOR2X1_19/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6001 XNOR2X1_19/a_12_41# AND2X2_16/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6002 gnd XNOR2X1_19/A XNOR2X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6003 XNOR2X1_19/a_18_6# XNOR2X1_19/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6004 AOI22X1_35/A XNOR2X1_19/A XNOR2X1_19/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6005 XNOR2X1_19/a_35_6# XNOR2X1_19/a_2_6# AOI22X1_35/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6006 gnd AND2X2_16/Y XNOR2X1_19/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6007 XNOR2X1_19/a_12_41# AND2X2_16/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6008 AND2X2_16/a_2_6# XOR2X1_40/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6009 vdd NAND3X1_8/C AND2X2_16/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6010 AND2X2_16/Y AND2X2_16/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6011 AND2X2_16/a_9_6# XOR2X1_40/A AND2X2_16/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6012 gnd NAND3X1_8/C AND2X2_16/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6013 AND2X2_16/Y AND2X2_16/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6014 vdd XOR2X1_40/A XOR2X1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6015 XOR2X1_40/a_18_54# XOR2X1_40/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6016 XOR2X1_40/Y XOR2X1_40/A XOR2X1_40/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6017 XOR2X1_40/a_35_54# XOR2X1_40/a_2_6# XOR2X1_40/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6018 vdd NAND3X1_8/C XOR2X1_40/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6019 XOR2X1_40/a_13_43# NAND3X1_8/C vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6020 gnd XOR2X1_40/A XOR2X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6021 XOR2X1_40/a_18_6# XOR2X1_40/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6022 XOR2X1_40/Y XOR2X1_40/a_2_6# XOR2X1_40/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6023 XOR2X1_40/a_35_6# XOR2X1_40/A XOR2X1_40/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6024 gnd NAND3X1_8/C XOR2X1_40/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6025 XOR2X1_40/a_13_43# NAND3X1_8/C gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6026 vdd INVX2_50/Y XOR2X1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6027 XOR2X1_39/a_18_54# XOR2X1_39/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6028 XOR2X1_39/Y INVX2_50/Y XOR2X1_39/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6029 XOR2X1_39/a_35_54# XOR2X1_39/a_2_6# XOR2X1_39/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6030 vdd INVX2_28/Y XOR2X1_39/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6031 XOR2X1_39/a_13_43# INVX2_28/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6032 gnd INVX2_50/Y XOR2X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6033 XOR2X1_39/a_18_6# XOR2X1_39/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6034 XOR2X1_39/Y XOR2X1_39/a_2_6# XOR2X1_39/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6035 XOR2X1_39/a_35_6# INVX2_50/Y XOR2X1_39/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6036 gnd INVX2_28/Y XOR2X1_39/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6037 XOR2X1_39/a_13_43# INVX2_28/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6038 vdd XOR2X1_69/B XNOR2X1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6039 XNOR2X1_17/a_18_54# XNOR2X1_17/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6040 XOR2X1_28/B XNOR2X1_17/a_2_6# XNOR2X1_17/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6041 XNOR2X1_17/a_35_54# XOR2X1_69/B XOR2X1_28/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6042 vdd XOR2X1_39/Y XNOR2X1_17/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6043 XNOR2X1_17/a_12_41# XOR2X1_39/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6044 gnd XOR2X1_69/B XNOR2X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6045 XNOR2X1_17/a_18_6# XNOR2X1_17/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6046 XOR2X1_28/B XOR2X1_69/B XNOR2X1_17/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6047 XNOR2X1_17/a_35_6# XNOR2X1_17/a_2_6# XOR2X1_28/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6048 gnd XOR2X1_39/Y XNOR2X1_17/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6049 XNOR2X1_17/a_12_41# XOR2X1_39/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6050 vdd XOR2X1_39/Y AOI22X1_32/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6051 AOI22X1_32/a_2_54# out_MuxData[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6052 NOR2X1_8/B out_MuxData[13] AOI22X1_32/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6053 AOI22X1_32/a_2_54# out_MuxData[14] NOR2X1_8/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6054 AOI22X1_32/a_11_6# XOR2X1_39/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6055 NOR2X1_8/B out_MuxData[9] AOI22X1_32/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6056 AOI22X1_32/a_28_6# out_MuxData[13] NOR2X1_8/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6057 gnd out_MuxData[14] AOI22X1_32/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6058 vdd INVX2_106/Y AOI22X1_31/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6059 AOI22X1_31/a_2_54# XOR2X1_27/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6060 NAND3X1_14/A XOR2X1_29/Y AOI22X1_31/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6061 AOI22X1_31/a_2_54# INVX2_71/Y NAND3X1_14/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6062 AOI22X1_31/a_11_6# INVX2_106/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6063 NAND3X1_14/A XOR2X1_27/Y AOI22X1_31/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6064 AOI22X1_31/a_28_6# XOR2X1_29/Y NAND3X1_14/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6065 gnd INVX2_71/Y AOI22X1_31/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6066 vdd out_MuxData[5] XOR2X1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6067 XOR2X1_35/a_18_54# XOR2X1_35/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6068 XOR2X1_35/Y out_MuxData[5] XOR2X1_35/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6069 XOR2X1_35/a_35_54# XOR2X1_35/a_2_6# XOR2X1_35/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6070 vdd out_MuxData[11] XOR2X1_35/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6071 XOR2X1_35/a_13_43# out_MuxData[11] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6072 gnd out_MuxData[5] XOR2X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6073 XOR2X1_35/a_18_6# XOR2X1_35/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6074 XOR2X1_35/Y XOR2X1_35/a_2_6# XOR2X1_35/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6075 XOR2X1_35/a_35_6# out_MuxData[5] XOR2X1_35/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6076 gnd out_MuxData[11] XOR2X1_35/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6077 XOR2X1_35/a_13_43# out_MuxData[11] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6078 OAI21X1_32/C XOR2X1_33/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6079 vdd NAND2X1_13/Y OAI21X1_32/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6080 OAI21X1_32/C XOR2X1_33/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6081 NAND3X1_13/a_9_6# XOR2X1_33/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6082 NAND3X1_13/a_14_6# NAND2X1_13/Y NAND3X1_13/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6083 OAI21X1_32/C XOR2X1_33/B NAND3X1_13/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6084 NAND2X1_13/Y AOI22X1_41/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6085 vdd XNOR2X1_24/Y NAND2X1_13/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6086 NAND2X1_13/a_9_6# AOI22X1_41/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6087 NAND2X1_13/Y XNOR2X1_24/Y NAND2X1_13/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6088 AND2X2_15/a_2_6# XOR2X1_33/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6089 vdd XOR2X1_33/B AND2X2_15/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6090 AND2X2_15/Y AND2X2_15/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6091 AND2X2_15/a_9_6# XOR2X1_33/A AND2X2_15/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6092 gnd XOR2X1_33/B AND2X2_15/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6093 AND2X2_15/Y AND2X2_15/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6094 vdd XOR2X1_33/A XOR2X1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6095 XOR2X1_33/a_18_54# XOR2X1_33/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6096 XOR2X1_33/Y XOR2X1_33/A XOR2X1_33/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6097 XOR2X1_33/a_35_54# XOR2X1_33/a_2_6# XOR2X1_33/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6098 vdd XOR2X1_33/B XOR2X1_33/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6099 XOR2X1_33/a_13_43# XOR2X1_33/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6100 gnd XOR2X1_33/A XOR2X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6101 XOR2X1_33/a_18_6# XOR2X1_33/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6102 XOR2X1_33/Y XOR2X1_33/a_2_6# XOR2X1_33/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6103 XOR2X1_33/a_35_6# XOR2X1_33/A XOR2X1_33/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6104 gnd XOR2X1_33/B XOR2X1_33/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6105 XOR2X1_33/a_13_43# XOR2X1_33/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6106 vdd BUFX2_11/Y DFFPOSX1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6107 DFFPOSX1_23/a_17_74# OAI21X1_31/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6108 DFFPOSX1_23/a_22_6# BUFX2_11/Y DFFPOSX1_23/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6109 DFFPOSX1_23/a_31_74# DFFPOSX1_23/a_2_6# DFFPOSX1_23/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6110 vdd DFFPOSX1_23/a_34_4# DFFPOSX1_23/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6111 DFFPOSX1_23/a_34_4# DFFPOSX1_23/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6112 DFFPOSX1_23/a_61_74# DFFPOSX1_23/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6113 DFFPOSX1_23/a_66_6# DFFPOSX1_23/a_2_6# DFFPOSX1_23/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6114 DFFPOSX1_23/a_76_84# BUFX2_11/Y DFFPOSX1_23/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6115 vdd out_MemBData[3] DFFPOSX1_23/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6116 gnd BUFX2_11/Y DFFPOSX1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6117 out_MemBData[3] DFFPOSX1_23/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6118 DFFPOSX1_23/a_17_6# OAI21X1_31/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6119 DFFPOSX1_23/a_22_6# DFFPOSX1_23/a_2_6# DFFPOSX1_23/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6120 DFFPOSX1_23/a_31_6# BUFX2_11/Y DFFPOSX1_23/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6121 gnd DFFPOSX1_23/a_34_4# DFFPOSX1_23/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6122 DFFPOSX1_23/a_34_4# DFFPOSX1_23/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6123 DFFPOSX1_23/a_61_6# DFFPOSX1_23/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6124 DFFPOSX1_23/a_66_6# BUFX2_11/Y DFFPOSX1_23/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6125 DFFPOSX1_23/a_76_6# DFFPOSX1_23/a_2_6# DFFPOSX1_23/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6126 gnd out_MemBData[3] DFFPOSX1_23/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6127 out_MemBData[3] DFFPOSX1_23/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6128 OAI21X1_30/a_9_54# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6129 OAI21X1_30/Y OR2X2_0/Y OAI21X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6130 vdd OAI21X1_30/C OAI21X1_30/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6131 gnd INVX2_25/A OAI21X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6132 OAI21X1_30/a_2_6# OR2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6133 OAI21X1_30/Y OAI21X1_30/C OAI21X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6134 vdd in_clkb DFFPOSX1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6135 DFFPOSX1_18/a_17_74# OAI21X1_29/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6136 DFFPOSX1_18/a_22_6# in_clkb DFFPOSX1_18/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6137 DFFPOSX1_18/a_31_74# DFFPOSX1_18/a_2_6# DFFPOSX1_18/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6138 vdd DFFPOSX1_18/a_34_4# DFFPOSX1_18/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6139 DFFPOSX1_18/a_34_4# DFFPOSX1_18/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6140 DFFPOSX1_18/a_61_74# DFFPOSX1_18/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6141 DFFPOSX1_18/a_66_6# DFFPOSX1_18/a_2_6# DFFPOSX1_18/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6142 DFFPOSX1_18/a_76_84# in_clkb DFFPOSX1_18/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6143 vdd out_temp_addNum[2] DFFPOSX1_18/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6144 gnd in_clkb DFFPOSX1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6145 out_temp_addNum[2] DFFPOSX1_18/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6146 DFFPOSX1_18/a_17_6# OAI21X1_29/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6147 DFFPOSX1_18/a_22_6# DFFPOSX1_18/a_2_6# DFFPOSX1_18/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6148 DFFPOSX1_18/a_31_6# in_clkb DFFPOSX1_18/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6149 gnd DFFPOSX1_18/a_34_4# DFFPOSX1_18/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6150 DFFPOSX1_18/a_34_4# DFFPOSX1_18/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6151 DFFPOSX1_18/a_61_6# DFFPOSX1_18/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6152 DFFPOSX1_18/a_66_6# in_clkb DFFPOSX1_18/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6153 DFFPOSX1_18/a_76_6# DFFPOSX1_18/a_2_6# DFFPOSX1_18/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6154 gnd out_temp_addNum[2] DFFPOSX1_18/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6155 out_temp_addNum[2] DFFPOSX1_18/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6156 OAI21X1_29/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6157 OAI21X1_29/Y INVX2_44/A OAI21X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6158 vdd NAND2X1_10/Y OAI21X1_29/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6159 gnd con_restart OAI21X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6160 OAI21X1_29/a_2_6# INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6161 OAI21X1_29/Y NAND2X1_10/Y OAI21X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6162 NAND2X1_10/Y out_temp_addNum[2] vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6163 vdd con_restart NAND2X1_10/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6164 NAND2X1_10/a_9_6# out_temp_addNum[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6165 NAND2X1_10/Y con_restart NAND2X1_10/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6166 vdd INVX2_41/Y DFFPOSX1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6167 DFFPOSX1_17/a_17_74# INVX2_36/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6168 DFFPOSX1_17/a_22_6# INVX2_41/Y DFFPOSX1_17/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6169 DFFPOSX1_17/a_31_74# DFFPOSX1_17/a_2_6# DFFPOSX1_17/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6170 vdd DFFPOSX1_17/a_34_4# DFFPOSX1_17/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6171 DFFPOSX1_17/a_34_4# DFFPOSX1_17/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6172 DFFPOSX1_17/a_61_74# DFFPOSX1_17/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6173 DFFPOSX1_17/a_66_6# DFFPOSX1_17/a_2_6# DFFPOSX1_17/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6174 DFFPOSX1_17/a_76_84# INVX2_41/Y DFFPOSX1_17/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6175 vdd con_countWriteout[0] DFFPOSX1_17/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6176 gnd INVX2_41/Y DFFPOSX1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6177 con_countWriteout[0] DFFPOSX1_17/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6178 DFFPOSX1_17/a_17_6# INVX2_36/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6179 DFFPOSX1_17/a_22_6# DFFPOSX1_17/a_2_6# DFFPOSX1_17/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6180 DFFPOSX1_17/a_31_6# INVX2_41/Y DFFPOSX1_17/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6181 gnd DFFPOSX1_17/a_34_4# DFFPOSX1_17/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6182 DFFPOSX1_17/a_34_4# DFFPOSX1_17/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6183 DFFPOSX1_17/a_61_6# DFFPOSX1_17/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6184 DFFPOSX1_17/a_66_6# INVX2_41/Y DFFPOSX1_17/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6185 DFFPOSX1_17/a_76_6# DFFPOSX1_17/a_2_6# DFFPOSX1_17/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6186 gnd con_countWriteout[0] DFFPOSX1_17/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6187 con_countWriteout[0] DFFPOSX1_17/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6188 INVX2_36/Y INVX2_36/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6189 INVX2_36/Y INVX2_36/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6190 vdd con_countWriteout[0] AOI22X1_29/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6191 AOI22X1_29/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6192 INVX2_36/A INVX2_11/A AOI22X1_29/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6193 AOI22X1_29/a_2_54# AOI22X1_29/C INVX2_36/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6194 AOI22X1_29/a_11_6# con_countWriteout[0] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6195 INVX2_36/A INVX2_11/Y AOI22X1_29/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6196 AOI22X1_29/a_28_6# INVX2_11/A INVX2_36/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6197 gnd AOI22X1_29/C AOI22X1_29/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6198 vdd BUFX2_9/Y DFFPOSX1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6199 DFFPOSX1_16/a_17_74# AND2X2_10/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6200 DFFPOSX1_16/a_22_6# BUFX2_9/Y DFFPOSX1_16/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6201 DFFPOSX1_16/a_31_74# DFFPOSX1_16/a_2_6# DFFPOSX1_16/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6202 vdd DFFPOSX1_16/a_34_4# DFFPOSX1_16/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6203 DFFPOSX1_16/a_34_4# DFFPOSX1_16/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6204 DFFPOSX1_16/a_61_74# DFFPOSX1_16/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6205 DFFPOSX1_16/a_66_6# DFFPOSX1_16/a_2_6# DFFPOSX1_16/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6206 DFFPOSX1_16/a_76_84# BUFX2_9/Y DFFPOSX1_16/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6207 vdd AOI22X1_29/C DFFPOSX1_16/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6208 gnd BUFX2_9/Y DFFPOSX1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6209 AOI22X1_29/C DFFPOSX1_16/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6210 DFFPOSX1_16/a_17_6# AND2X2_10/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6211 DFFPOSX1_16/a_22_6# DFFPOSX1_16/a_2_6# DFFPOSX1_16/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6212 DFFPOSX1_16/a_31_6# BUFX2_9/Y DFFPOSX1_16/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6213 gnd DFFPOSX1_16/a_34_4# DFFPOSX1_16/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6214 DFFPOSX1_16/a_34_4# DFFPOSX1_16/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6215 DFFPOSX1_16/a_61_6# DFFPOSX1_16/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6216 DFFPOSX1_16/a_66_6# BUFX2_9/Y DFFPOSX1_16/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6217 DFFPOSX1_16/a_76_6# DFFPOSX1_16/a_2_6# DFFPOSX1_16/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6218 gnd AOI22X1_29/C DFFPOSX1_16/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6219 AOI22X1_29/C DFFPOSX1_16/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6220 OAI21X1_28/a_9_54# OAI21X1_28/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6221 INVX2_35/A INVX2_22/Y OAI21X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6222 vdd AOI21X1_3/Y INVX2_35/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6223 gnd OAI21X1_28/A OAI21X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6224 OAI21X1_28/a_2_6# INVX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6225 INVX2_35/A AOI21X1_3/Y OAI21X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6226 AND2X2_6/B in_reset vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6227 AND2X2_6/B in_reset gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6228 vdd NOR2X1_5/Y AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M6229 AOI21X1_3/a_2_54# in_inp vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6230 AOI21X1_3/Y in_reset AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6231 AOI21X1_3/a_12_6# NOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6232 AOI21X1_3/Y in_inp AOI21X1_3/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M6233 gnd in_reset AOI21X1_3/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6234 INVX2_21/A INVX2_32/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6235 vdd INVX2_34/Y INVX2_21/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6236 INVX2_21/A INVX2_31/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6237 NAND3X1_11/a_9_6# INVX2_32/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6238 NAND3X1_11/a_14_6# INVX2_34/Y NAND3X1_11/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6239 INVX2_21/A INVX2_31/Y NAND3X1_11/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6240 OAI21X1_28/A out_state[0] vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6241 vdd INVX2_32/Y OAI21X1_28/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6242 OAI21X1_28/A out_state[2] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6243 NAND3X1_10/a_9_6# out_state[0] gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6244 NAND3X1_10/a_14_6# INVX2_32/Y NAND3X1_10/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6245 OAI21X1_28/A out_state[2] NAND3X1_10/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6246 INVX2_32/Y out_state[1] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6247 INVX2_32/Y out_state[1] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6248 INVX2_19/A out_state[2] vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6249 vdd INVX2_31/Y INVX2_19/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6250 INVX2_19/A out_state[1] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6251 NAND3X1_9/a_9_6# out_state[2] gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6252 NAND3X1_9/a_14_6# INVX2_31/Y NAND3X1_9/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6253 INVX2_19/A out_state[1] NAND3X1_9/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6254 INVX2_31/Y out_state[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6255 INVX2_31/Y out_state[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6256 NAND2X1_9/Y NAND2X1_9/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6257 vdd AOI21X1_4/Y NAND2X1_9/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6258 NAND2X1_9/a_9_6# NAND2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6259 NAND2X1_9/Y AOI21X1_4/Y NAND2X1_9/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6260 vdd out_MuxData[5] XOR2X1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6261 XOR2X1_32/a_18_54# XOR2X1_32/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6262 XOR2X1_32/Y out_MuxData[5] XOR2X1_32/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6263 XOR2X1_32/a_35_54# XOR2X1_32/a_2_6# XOR2X1_32/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6264 vdd out_MuxData[6] XOR2X1_32/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6265 XOR2X1_32/a_13_43# out_MuxData[6] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6266 gnd out_MuxData[5] XOR2X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6267 XOR2X1_32/a_18_6# XOR2X1_32/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6268 XOR2X1_32/Y XOR2X1_32/a_2_6# XOR2X1_32/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6269 XOR2X1_32/a_35_6# out_MuxData[5] XOR2X1_32/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6270 gnd out_MuxData[6] XOR2X1_32/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6271 XOR2X1_32/a_13_43# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6272 NAND2X1_8/Y out_MuxData[5] vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6273 vdd out_MuxData[4] NAND2X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6274 NAND2X1_8/a_9_6# out_MuxData[5] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6275 NAND2X1_8/Y out_MuxData[4] NAND2X1_8/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6276 OAI21X1_26/a_9_54# XOR2X1_81/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6277 INVX2_29/A XNOR2X1_22/A OAI21X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6278 vdd NAND2X1_8/Y INVX2_29/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6279 gnd XOR2X1_81/A OAI21X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6280 OAI21X1_26/a_2_6# XNOR2X1_22/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6281 INVX2_29/A NAND2X1_8/Y OAI21X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6282 vdd XOR2X1_81/A XNOR2X1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6283 XNOR2X1_16/a_18_54# XNOR2X1_16/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6284 XOR2X1_43/B XNOR2X1_16/a_2_6# XNOR2X1_16/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6285 XNOR2X1_16/a_35_54# XOR2X1_81/A XOR2X1_43/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6286 vdd XOR2X1_32/Y XNOR2X1_16/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6287 XNOR2X1_16/a_12_41# XOR2X1_32/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6288 gnd XOR2X1_81/A XNOR2X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6289 XNOR2X1_16/a_18_6# XNOR2X1_16/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6290 XOR2X1_43/B XOR2X1_81/A XNOR2X1_16/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6291 XNOR2X1_16/a_35_6# XNOR2X1_16/a_2_6# XOR2X1_43/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6292 gnd XOR2X1_32/Y XNOR2X1_16/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6293 XNOR2X1_16/a_12_41# XOR2X1_32/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6294 vdd XOR2X1_43/B AOI22X1_28/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6295 AOI22X1_28/a_2_54# out_MuxData[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6296 NOR2X1_12/A out_MuxData[14] AOI22X1_28/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6297 AOI22X1_28/a_2_54# XOR2X1_43/Y NOR2X1_12/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6298 AOI22X1_28/a_11_6# XOR2X1_43/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6299 NOR2X1_12/A out_MuxData[15] AOI22X1_28/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6300 AOI22X1_28/a_28_6# out_MuxData[14] NOR2X1_12/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6301 gnd XOR2X1_43/Y AOI22X1_28/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6302 NOR2X1_9/A INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6303 NOR2X1_9/A INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6304 vdd INVX2_29/A XOR2X1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6305 XOR2X1_31/a_18_54# XOR2X1_31/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6306 NAND2X1_7/A INVX2_29/A XOR2X1_31/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6307 XOR2X1_31/a_35_54# XOR2X1_31/a_2_6# NAND2X1_7/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6308 vdd NOR2X1_9/B XOR2X1_31/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6309 XOR2X1_31/a_13_43# NOR2X1_9/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6310 gnd INVX2_29/A XOR2X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6311 XOR2X1_31/a_18_6# XOR2X1_31/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6312 NAND2X1_7/A XOR2X1_31/a_2_6# XOR2X1_31/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6313 XOR2X1_31/a_35_6# INVX2_29/A NAND2X1_7/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6314 gnd NOR2X1_9/B XOR2X1_31/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6315 XOR2X1_31/a_13_43# NOR2X1_9/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6316 NOR2X1_9/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6317 NOR2X1_9/Y NOR2X1_9/B NOR2X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6318 NOR2X1_9/Y NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6319 gnd NOR2X1_9/B NOR2X1_9/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6320 vdd XOR2X1_29/A XOR2X1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6321 XOR2X1_29/a_18_54# XOR2X1_29/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6322 XOR2X1_29/Y XOR2X1_29/A XOR2X1_29/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6323 XOR2X1_29/a_35_54# XOR2X1_29/a_2_6# XOR2X1_29/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6324 vdd NOR2X1_9/Y XOR2X1_29/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6325 XOR2X1_29/a_13_43# NOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6326 gnd XOR2X1_29/A XOR2X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6327 XOR2X1_29/a_18_6# XOR2X1_29/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6328 XOR2X1_29/Y XOR2X1_29/a_2_6# XOR2X1_29/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6329 XOR2X1_29/a_35_6# XOR2X1_29/A XOR2X1_29/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6330 gnd NOR2X1_9/Y XOR2X1_29/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6331 XOR2X1_29/a_13_43# NOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6332 OAI21X1_23/a_9_54# INVX2_27/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6333 XOR2X1_29/A NAND2X1_7/A OAI21X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6334 vdd NAND3X1_8/Y XOR2X1_29/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6335 gnd INVX2_27/Y OAI21X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6336 OAI21X1_23/a_2_6# NAND2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6337 XOR2X1_29/A NAND3X1_8/Y OAI21X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6338 OAI21X1_22/a_9_54# INVX2_27/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6339 XNOR2X1_19/A NAND2X1_7/A OAI21X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6340 vdd NAND3X1_8/B XNOR2X1_19/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6341 gnd INVX2_27/Y OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6342 OAI21X1_22/a_2_6# NAND2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6343 XNOR2X1_19/A NAND3X1_8/B OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6344 NAND3X1_8/Y XOR2X1_40/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6345 vdd NAND3X1_8/B NAND3X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6346 NAND3X1_8/Y NAND3X1_8/C vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6347 NAND3X1_8/a_9_6# XOR2X1_40/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6348 NAND3X1_8/a_14_6# NAND3X1_8/B NAND3X1_8/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6349 NAND3X1_8/Y NAND3X1_8/C NAND3X1_8/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6350 vdd XNOR2X1_9/A XNOR2X1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6351 XNOR2X1_14/a_18_54# XNOR2X1_14/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6352 NAND3X1_8/C XNOR2X1_14/a_2_6# XNOR2X1_14/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6353 XNOR2X1_14/a_35_54# XNOR2X1_9/A NAND3X1_8/C vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6354 vdd INVX2_39/A XNOR2X1_14/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6355 XNOR2X1_14/a_12_41# INVX2_39/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6356 gnd XNOR2X1_9/A XNOR2X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6357 XNOR2X1_14/a_18_6# XNOR2X1_14/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6358 NAND3X1_8/C XNOR2X1_9/A XNOR2X1_14/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6359 XNOR2X1_14/a_35_6# XNOR2X1_14/a_2_6# NAND3X1_8/C Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6360 gnd INVX2_39/A XNOR2X1_14/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6361 XNOR2X1_14/a_12_41# INVX2_39/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6362 vdd XOR2X1_28/B AOI22X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6363 AOI22X1_25/a_2_54# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6364 NOR2X1_8/A out_MuxData[6] AOI22X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6365 AOI22X1_25/a_2_54# XOR2X1_28/Y NOR2X1_8/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6366 AOI22X1_25/a_11_6# XOR2X1_28/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6367 NOR2X1_8/A out_MuxData[7] AOI22X1_25/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6368 AOI22X1_25/a_28_6# out_MuxData[6] NOR2X1_8/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6369 gnd XOR2X1_28/Y AOI22X1_25/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6370 NOR2X1_8/a_9_54# NOR2X1_8/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6371 NOR2X1_8/Y NOR2X1_8/B NOR2X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6372 NOR2X1_8/Y NOR2X1_8/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6373 gnd NOR2X1_8/B NOR2X1_8/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6374 vdd XOR2X1_27/A XOR2X1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6375 XOR2X1_27/a_18_54# XOR2X1_27/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6376 XOR2X1_27/Y XOR2X1_27/A XOR2X1_27/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6377 XOR2X1_27/a_35_54# XOR2X1_27/a_2_6# XOR2X1_27/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6378 vdd NOR2X1_8/Y XOR2X1_27/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6379 XOR2X1_27/a_13_43# NOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6380 gnd XOR2X1_27/A XOR2X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6381 XOR2X1_27/a_18_6# XOR2X1_27/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6382 XOR2X1_27/Y XOR2X1_27/a_2_6# XOR2X1_27/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6383 XOR2X1_27/a_35_6# XOR2X1_27/A XOR2X1_27/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6384 gnd NOR2X1_8/Y XOR2X1_27/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6385 XOR2X1_27/a_13_43# NOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6386 OAI21X1_21/a_9_54# AOI22X1_41/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6387 XNOR2X1_11/A XNOR2X1_24/Y OAI21X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6388 vdd NAND2X1_13/Y XNOR2X1_11/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6389 gnd AOI22X1_41/Y OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6390 OAI21X1_21/a_2_6# XNOR2X1_24/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6391 XNOR2X1_11/A NAND2X1_13/Y OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6392 vdd XNOR2X1_11/A XNOR2X1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6393 XNOR2X1_11/a_18_54# XNOR2X1_11/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6394 AOI22X1_23/A XNOR2X1_11/a_2_6# XNOR2X1_11/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6395 XNOR2X1_11/a_35_54# XNOR2X1_11/A AOI22X1_23/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6396 vdd AND2X2_15/Y XNOR2X1_11/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6397 XNOR2X1_11/a_12_41# AND2X2_15/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6398 gnd XNOR2X1_11/A XNOR2X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6399 XNOR2X1_11/a_18_6# XNOR2X1_11/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6400 AOI22X1_23/A XNOR2X1_11/A XNOR2X1_11/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6401 XNOR2X1_11/a_35_6# XNOR2X1_11/a_2_6# AOI22X1_23/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6402 gnd AND2X2_15/Y XNOR2X1_11/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6403 XNOR2X1_11/a_12_41# AND2X2_15/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6404 vdd AOI22X1_23/A AOI22X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6405 AOI22X1_23/a_2_54# INVX2_104/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6406 AND2X2_13/A INVX2_93/Y AOI22X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6407 AOI22X1_23/a_2_54# XNOR2X1_0/Y AND2X2_13/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6408 AOI22X1_23/a_11_6# AOI22X1_23/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6409 AND2X2_13/A INVX2_104/Y AOI22X1_23/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6410 AOI22X1_23/a_28_6# INVX2_93/Y AND2X2_13/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6411 gnd XNOR2X1_0/Y AOI22X1_23/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6412 vdd INVX2_93/Y AOI22X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6413 AOI22X1_22/a_2_54# XOR2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6414 NAND3X1_7/B XOR2X1_33/Y AOI22X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6415 AOI22X1_22/a_2_54# INVX2_104/Y NAND3X1_7/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6416 AOI22X1_22/a_11_6# INVX2_93/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6417 NAND3X1_7/B XOR2X1_1/Y AOI22X1_22/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6418 AOI22X1_22/a_28_6# XOR2X1_33/Y NAND3X1_7/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6419 gnd INVX2_104/Y AOI22X1_22/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6420 NAND3X1_7/Y NAND3X1_7/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6421 vdd NAND3X1_7/B NAND3X1_7/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6422 NAND3X1_7/Y AND2X2_21/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6423 NAND3X1_7/a_9_6# NAND3X1_7/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6424 NAND3X1_7/a_14_6# NAND3X1_7/B NAND3X1_7/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6425 NAND3X1_7/Y AND2X2_21/Y NAND3X1_7/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6426 OAI21X1_20/a_9_54# NOR2X1_7/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6427 OAI21X1_31/C AND2X2_19/Y OAI21X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6428 vdd out_MemBData[3] OAI21X1_31/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6429 gnd NOR2X1_7/Y OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6430 OAI21X1_20/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6431 OAI21X1_31/C out_MemBData[3] OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6432 NOR2X1_6/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6433 NOR2X1_6/Y INVX2_25/Y NOR2X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6434 NOR2X1_6/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6435 gnd INVX2_25/Y NOR2X1_6/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6436 OAI21X1_19/a_9_54# NOR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6437 OAI21X1_30/C AND2X2_19/Y OAI21X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6438 vdd out_MemBData[1] OAI21X1_30/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6439 gnd NOR2X1_6/Y OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6440 OAI21X1_19/a_2_6# AND2X2_19/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6441 OAI21X1_30/C out_MemBData[1] OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6442 INVX2_25/Y INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6443 INVX2_25/Y INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6444 vdd BUFX2_9/Y DFFPOSX1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6445 DFFPOSX1_15/a_17_74# AND2X2_11/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6446 DFFPOSX1_15/a_22_6# BUFX2_9/Y DFFPOSX1_15/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6447 DFFPOSX1_15/a_31_74# DFFPOSX1_15/a_2_6# DFFPOSX1_15/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6448 vdd DFFPOSX1_15/a_34_4# DFFPOSX1_15/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6449 DFFPOSX1_15/a_34_4# DFFPOSX1_15/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6450 DFFPOSX1_15/a_61_74# DFFPOSX1_15/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6451 DFFPOSX1_15/a_66_6# DFFPOSX1_15/a_2_6# DFFPOSX1_15/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6452 DFFPOSX1_15/a_76_84# BUFX2_9/Y DFFPOSX1_15/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6453 vdd AOI22X1_19/C DFFPOSX1_15/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6454 gnd BUFX2_9/Y DFFPOSX1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6455 AOI22X1_19/C DFFPOSX1_15/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6456 DFFPOSX1_15/a_17_6# AND2X2_11/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6457 DFFPOSX1_15/a_22_6# DFFPOSX1_15/a_2_6# DFFPOSX1_15/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6458 DFFPOSX1_15/a_31_6# BUFX2_9/Y DFFPOSX1_15/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6459 gnd DFFPOSX1_15/a_34_4# DFFPOSX1_15/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6460 DFFPOSX1_15/a_34_4# DFFPOSX1_15/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6461 DFFPOSX1_15/a_61_6# DFFPOSX1_15/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6462 DFFPOSX1_15/a_66_6# BUFX2_9/Y DFFPOSX1_15/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6463 DFFPOSX1_15/a_76_6# DFFPOSX1_15/a_2_6# DFFPOSX1_15/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6464 gnd AOI22X1_19/C DFFPOSX1_15/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6465 AOI22X1_19/C DFFPOSX1_15/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6466 AND2X2_12/a_2_6# HAX1_5/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6467 vdd AND2X2_6/B AND2X2_12/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6468 AND2X2_12/Y AND2X2_12/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6469 AND2X2_12/a_9_6# HAX1_5/YS AND2X2_12/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6470 gnd AND2X2_6/B AND2X2_12/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6471 AND2X2_12/Y AND2X2_12/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6472 vdd BUFX2_9/Y DFFPOSX1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6473 DFFPOSX1_14/a_17_74# AND2X2_12/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6474 DFFPOSX1_14/a_22_6# BUFX2_9/Y DFFPOSX1_14/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6475 DFFPOSX1_14/a_31_74# DFFPOSX1_14/a_2_6# DFFPOSX1_14/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6476 vdd DFFPOSX1_14/a_34_4# DFFPOSX1_14/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6477 DFFPOSX1_14/a_34_4# DFFPOSX1_14/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6478 DFFPOSX1_14/a_61_74# DFFPOSX1_14/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6479 DFFPOSX1_14/a_66_6# DFFPOSX1_14/a_2_6# DFFPOSX1_14/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6480 DFFPOSX1_14/a_76_84# BUFX2_9/Y DFFPOSX1_14/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6481 vdd AOI22X1_18/C DFFPOSX1_14/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6482 gnd BUFX2_9/Y DFFPOSX1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6483 AOI22X1_18/C DFFPOSX1_14/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6484 DFFPOSX1_14/a_17_6# AND2X2_12/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6485 DFFPOSX1_14/a_22_6# DFFPOSX1_14/a_2_6# DFFPOSX1_14/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6486 DFFPOSX1_14/a_31_6# BUFX2_9/Y DFFPOSX1_14/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6487 gnd DFFPOSX1_14/a_34_4# DFFPOSX1_14/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6488 DFFPOSX1_14/a_34_4# DFFPOSX1_14/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6489 DFFPOSX1_14/a_61_6# DFFPOSX1_14/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6490 DFFPOSX1_14/a_66_6# BUFX2_9/Y DFFPOSX1_14/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6491 DFFPOSX1_14/a_76_6# DFFPOSX1_14/a_2_6# DFFPOSX1_14/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6492 gnd AOI22X1_18/C DFFPOSX1_14/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6493 AOI22X1_18/C DFFPOSX1_14/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6494 INVX2_22/Y con_loseSig vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6495 INVX2_22/Y con_loseSig gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6496 OAI21X1_17/a_9_54# OAI21X1_28/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6497 AOI21X1_4/C OAI21X1_18/Y OAI21X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6498 vdd AND2X2_6/B AOI21X1_4/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6499 gnd OAI21X1_28/A OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6500 OAI21X1_17/a_2_6# OAI21X1_18/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6501 AOI21X1_4/C AND2X2_6/B OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6502 NOR2X1_5/a_9_54# out_state[2] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6503 NOR2X1_5/Y out_state[1] NOR2X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6504 NOR2X1_5/Y out_state[2] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6505 gnd out_state[1] NOR2X1_5/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6506 INVX2_21/Y INVX2_21/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6507 INVX2_21/Y INVX2_21/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6508 INVX2_20/Y in_inp vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6509 INVX2_20/Y in_inp gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6510 INVX2_19/Y INVX2_19/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6511 INVX2_19/Y INVX2_19/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6512 vdd INVX2_21/Y AOI22X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6513 AOI22X1_17/a_2_54# NAND3X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6514 NAND2X1_9/A INVX2_19/Y AOI22X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6515 AOI22X1_17/a_2_54# in_inp NAND2X1_9/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6516 AOI22X1_17/a_11_6# INVX2_21/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6517 NAND2X1_9/A NAND3X1_5/Y AOI22X1_17/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6518 AOI22X1_17/a_28_6# INVX2_19/Y NAND2X1_9/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6519 gnd in_inp AOI22X1_17/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6520 INVX2_30/Y INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6521 INVX2_30/Y INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6522 OAI21X1_25/a_9_54# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6523 XNOR2X1_22/A out_MuxData[4] OAI21X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6524 vdd NAND2X1_8/Y XNOR2X1_22/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6525 gnd out_MuxData[5] OAI21X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6526 OAI21X1_25/a_2_6# out_MuxData[4] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6527 XNOR2X1_22/A NAND2X1_8/Y OAI21X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6528 OAI21X1_24/a_9_54# OAI22X1_6/C vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6529 INVX2_30/A XNOR2X1_22/A OAI21X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6530 vdd NAND2X1_8/Y INVX2_30/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6531 gnd OAI22X1_6/C OAI21X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6532 OAI21X1_24/a_2_6# XNOR2X1_22/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6533 INVX2_30/A NAND2X1_8/Y OAI21X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6534 vdd XNOR2X1_22/A XNOR2X1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6535 XNOR2X1_15/a_18_54# XNOR2X1_15/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6536 XOR2X1_23/A XNOR2X1_15/a_2_6# XNOR2X1_15/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6537 XNOR2X1_15/a_35_54# XNOR2X1_22/A XOR2X1_23/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6538 vdd out_MuxData[0] XNOR2X1_15/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6539 XNOR2X1_15/a_12_41# out_MuxData[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6540 gnd XNOR2X1_22/A XNOR2X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6541 XNOR2X1_15/a_18_6# XNOR2X1_15/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6542 XOR2X1_23/A XNOR2X1_22/A XNOR2X1_15/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6543 XNOR2X1_15/a_35_6# XNOR2X1_15/a_2_6# XOR2X1_23/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6544 gnd out_MuxData[0] XNOR2X1_15/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6545 XNOR2X1_15/a_12_41# out_MuxData[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6546 vdd out_MuxData[0] AOI22X1_27/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6547 AOI22X1_27/a_2_54# out_MuxData[14] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6548 OAI21X1_4/A out_MuxData[4] AOI22X1_27/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6549 AOI22X1_27/a_2_54# XOR2X1_30/Y OAI21X1_4/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6550 AOI22X1_27/a_11_6# out_MuxData[0] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6551 OAI21X1_4/A out_MuxData[14] AOI22X1_27/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6552 AOI22X1_27/a_28_6# out_MuxData[4] OAI21X1_4/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6553 gnd XOR2X1_30/Y AOI22X1_27/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6554 vdd OAI22X1_6/C XOR2X1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6555 XOR2X1_30/a_18_54# XOR2X1_30/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6556 XOR2X1_30/Y OAI22X1_6/C XOR2X1_30/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6557 XOR2X1_30/a_35_54# XOR2X1_30/a_2_6# XOR2X1_30/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6558 vdd INVX2_28/Y XOR2X1_30/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6559 XOR2X1_30/a_13_43# INVX2_28/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6560 gnd OAI22X1_6/C XOR2X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6561 XOR2X1_30/a_18_6# XOR2X1_30/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6562 XOR2X1_30/Y XOR2X1_30/a_2_6# XOR2X1_30/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6563 XOR2X1_30/a_35_6# OAI22X1_6/C XOR2X1_30/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6564 gnd INVX2_28/Y XOR2X1_30/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6565 XOR2X1_30/a_13_43# INVX2_28/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6566 INVX2_28/Y out_MuxData[14] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6567 INVX2_28/Y out_MuxData[14] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6568 vdd INVX2_25/Y AOI22X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6569 AOI22X1_26/a_2_54# XOR2X1_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6570 NAND3X1_17/B XOR2X1_7/Y AOI22X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6571 AOI22X1_26/a_2_54# INVX2_26/Y NAND3X1_17/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6572 AOI22X1_26/a_11_6# INVX2_25/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6573 NAND3X1_17/B XOR2X1_24/Y AOI22X1_26/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6574 AOI22X1_26/a_28_6# XOR2X1_7/Y NAND3X1_17/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6575 gnd INVX2_26/Y AOI22X1_26/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6576 NAND3X1_8/B NAND2X1_7/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6577 vdd INVX2_27/Y NAND3X1_8/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6578 NAND2X1_7/a_9_6# NAND2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6579 NAND3X1_8/B INVX2_27/Y NAND2X1_7/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6580 INVX2_27/Y INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6581 INVX2_27/Y INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6582 vdd out_MuxData[7] XOR2X1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6583 XOR2X1_28/a_18_54# XOR2X1_28/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6584 XOR2X1_28/Y out_MuxData[7] XOR2X1_28/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6585 XOR2X1_28/a_35_54# XOR2X1_28/a_2_6# XOR2X1_28/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6586 vdd XOR2X1_28/B XOR2X1_28/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6587 XOR2X1_28/a_13_43# XOR2X1_28/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6588 gnd out_MuxData[7] XOR2X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6589 XOR2X1_28/a_18_6# XOR2X1_28/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6590 XOR2X1_28/Y XOR2X1_28/a_2_6# XOR2X1_28/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6591 XOR2X1_28/a_35_6# out_MuxData[7] XOR2X1_28/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6592 gnd XOR2X1_28/B XOR2X1_28/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6593 XOR2X1_28/a_13_43# XOR2X1_28/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6594 vdd INVX2_16/Y XNOR2X1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6595 XNOR2X1_13/a_18_54# XNOR2X1_13/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6596 AND2X2_14/A XNOR2X1_13/a_2_6# XNOR2X1_13/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6597 XNOR2X1_13/a_35_54# INVX2_16/Y AND2X2_14/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6598 vdd XOR2X1_28/Y XNOR2X1_13/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6599 XNOR2X1_13/a_12_41# XOR2X1_28/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6600 gnd INVX2_16/Y XNOR2X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6601 XNOR2X1_13/a_18_6# XNOR2X1_13/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6602 AND2X2_14/A INVX2_16/Y XNOR2X1_13/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6603 XNOR2X1_13/a_35_6# XNOR2X1_13/a_2_6# AND2X2_14/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6604 gnd XOR2X1_28/Y XNOR2X1_13/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6605 XNOR2X1_13/a_12_41# XOR2X1_28/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6606 vdd out_MuxData[11] AOI22X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6607 AOI22X1_24/a_2_54# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6608 NAND2X1_4/A out_MuxData[15] AOI22X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6609 AOI22X1_24/a_2_54# XOR2X1_35/Y NAND2X1_4/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6610 AOI22X1_24/a_11_6# out_MuxData[11] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6611 NAND2X1_4/A out_MuxData[5] AOI22X1_24/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6612 AOI22X1_24/a_28_6# out_MuxData[15] NAND2X1_4/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6613 gnd XOR2X1_35/Y AOI22X1_24/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6614 vdd INVX2_5/A XNOR2X1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6615 XNOR2X1_12/a_18_54# XNOR2X1_12/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6616 NAND3X1_3/C XNOR2X1_12/a_2_6# XNOR2X1_12/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6617 XNOR2X1_12/a_35_54# INVX2_5/A NAND3X1_3/C vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6618 vdd XOR2X1_35/Y XNOR2X1_12/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6619 XNOR2X1_12/a_12_41# XOR2X1_35/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6620 gnd INVX2_5/A XNOR2X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6621 XNOR2X1_12/a_18_6# XNOR2X1_12/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6622 NAND3X1_3/C INVX2_5/A XNOR2X1_12/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6623 XNOR2X1_12/a_35_6# XNOR2X1_12/a_2_6# NAND3X1_3/C Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6624 gnd XOR2X1_35/Y XNOR2X1_12/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6625 XNOR2X1_12/a_12_41# XOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6626 vdd NAND3X1_3/C XOR2X1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6627 XOR2X1_26/a_18_54# XOR2X1_26/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6628 XOR2X1_26/Y NAND3X1_3/C XOR2X1_26/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6629 XOR2X1_26/a_35_54# XOR2X1_26/a_2_6# XOR2X1_26/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6630 vdd AND2X2_14/A XOR2X1_26/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6631 XOR2X1_26/a_13_43# AND2X2_14/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6632 gnd NAND3X1_3/C XOR2X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6633 XOR2X1_26/a_18_6# XOR2X1_26/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6634 XOR2X1_26/Y XOR2X1_26/a_2_6# XOR2X1_26/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6635 XOR2X1_26/a_35_6# NAND3X1_3/C XOR2X1_26/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6636 gnd AND2X2_14/A XOR2X1_26/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6637 XOR2X1_26/a_13_43# AND2X2_14/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6638 AND2X2_14/a_2_6# AND2X2_14/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6639 vdd NAND3X1_3/C AND2X2_14/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6640 AND2X2_14/Y AND2X2_14/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6641 AND2X2_14/a_9_6# AND2X2_14/A AND2X2_14/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6642 gnd NAND3X1_3/C AND2X2_14/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6643 AND2X2_14/Y AND2X2_14/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6644 AND2X2_13/a_2_6# AND2X2_13/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6645 vdd AND2X2_13/B AND2X2_13/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6646 AND2X2_13/Y AND2X2_13/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6647 AND2X2_13/a_9_6# AND2X2_13/A AND2X2_13/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6648 gnd AND2X2_13/B AND2X2_13/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6649 AND2X2_13/Y AND2X2_13/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6650 vdd XNOR2X1_8/Y AOI22X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6651 AOI22X1_21/a_2_54# INVX2_106/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6652 AND2X2_13/B NOR2X1_41/B AOI22X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6653 AOI22X1_21/a_2_54# XNOR2X1_7/Y AND2X2_13/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6654 AOI22X1_21/a_11_6# XNOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6655 AND2X2_13/B INVX2_106/Y AOI22X1_21/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6656 AOI22X1_21/a_28_6# NOR2X1_41/B AND2X2_13/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6657 gnd XNOR2X1_7/Y AOI22X1_21/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6658 vdd NOR2X1_41/B AOI22X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6659 AOI22X1_20/a_2_54# XOR2X1_13/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6660 NAND3X1_7/A XOR2X1_26/Y AOI22X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6661 AOI22X1_20/a_2_54# INVX2_106/Y NAND3X1_7/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6662 AOI22X1_20/a_11_6# NOR2X1_41/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6663 NAND3X1_7/A XOR2X1_13/Y AOI22X1_20/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6664 AOI22X1_20/a_28_6# XOR2X1_26/Y NAND3X1_7/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6665 gnd INVX2_106/Y AOI22X1_20/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6666 NOR2X1_7/a_9_54# con_restart vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6667 NOR2X1_7/Y INVX2_26/Y NOR2X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6668 NOR2X1_7/Y con_restart gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6669 gnd INVX2_26/Y NOR2X1_7/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6670 INVX2_26/Y INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6671 INVX2_26/Y INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6672 INVX2_24/Y INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6673 INVX2_24/Y INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6674 vdd con_countWriteout[2] AOI22X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6675 AOI22X1_19/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6676 INVX2_24/A INVX2_11/A AOI22X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6677 AOI22X1_19/a_2_54# AOI22X1_19/C INVX2_24/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6678 AOI22X1_19/a_11_6# con_countWriteout[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6679 INVX2_24/A INVX2_11/Y AOI22X1_19/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6680 AOI22X1_19/a_28_6# INVX2_11/A INVX2_24/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6681 gnd AOI22X1_19/C AOI22X1_19/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6682 AND2X2_11/a_2_6# HAX1_6/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6683 vdd AND2X2_6/B AND2X2_11/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6684 AND2X2_11/Y AND2X2_11/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6685 AND2X2_11/a_9_6# HAX1_6/YS AND2X2_11/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6686 gnd AND2X2_6/B AND2X2_11/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6687 AND2X2_11/Y AND2X2_11/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6688 vdd con_countWriteout[2] HAX1_6/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M6689 HAX1_6/a_2_74# HAX1_6/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6690 vdd HAX1_6/a_2_74# HAX1_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6691 HAX1_6/a_41_74# HAX1_6/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M6692 HAX1_6/a_49_54# HAX1_6/B HAX1_6/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6693 vdd con_countWriteout[2] HAX1_6/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6694 HAX1_6/YS HAX1_6/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6695 HAX1_6/a_9_6# con_countWriteout[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6696 HAX1_6/a_2_74# HAX1_6/B HAX1_6/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6697 gnd HAX1_6/a_2_74# HAX1_4/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M6698 HAX1_6/a_38_6# HAX1_6/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M6699 HAX1_6/a_41_74# HAX1_6/B HAX1_6/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6700 HAX1_6/a_38_6# con_countWriteout[2] HAX1_6/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6701 HAX1_6/YS HAX1_6/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6702 vdd con_countWriteout[1] HAX1_5/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M6703 HAX1_5/a_2_74# con_countWriteout[0] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6704 vdd HAX1_5/a_2_74# HAX1_6/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6705 HAX1_5/a_41_74# HAX1_5/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M6706 HAX1_5/a_49_54# con_countWriteout[0] HAX1_5/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6707 vdd con_countWriteout[1] HAX1_5/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6708 HAX1_5/YS HAX1_5/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6709 HAX1_5/a_9_6# con_countWriteout[1] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6710 HAX1_5/a_2_74# con_countWriteout[0] HAX1_5/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6711 gnd HAX1_5/a_2_74# HAX1_6/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M6712 HAX1_5/a_38_6# HAX1_5/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M6713 HAX1_5/a_41_74# con_countWriteout[0] HAX1_5/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6714 HAX1_5/a_38_6# con_countWriteout[1] HAX1_5/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6715 HAX1_5/YS HAX1_5/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6716 vdd con_countWriteout[1] AOI22X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6717 AOI22X1_18/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6718 INVX2_12/A INVX2_11/A AOI22X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6719 AOI22X1_18/a_2_54# AOI22X1_18/C INVX2_12/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6720 AOI22X1_18/a_11_6# con_countWriteout[1] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6721 INVX2_12/A INVX2_11/Y AOI22X1_18/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6722 AOI22X1_18/a_28_6# INVX2_11/A INVX2_12/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6723 gnd AOI22X1_18/C AOI22X1_18/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6724 INVX2_23/Y con_countWriteout[0] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6725 INVX2_23/Y con_countWriteout[0] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6726 AND2X2_10/a_2_6# INVX2_23/Y vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6727 vdd AND2X2_6/B AND2X2_10/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6728 AND2X2_10/Y AND2X2_10/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6729 AND2X2_10/a_9_6# INVX2_23/Y AND2X2_10/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6730 gnd AND2X2_6/B AND2X2_10/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6731 AND2X2_10/Y AND2X2_10/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6732 OAI21X1_18/a_9_54# INVX2_10/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6733 OAI21X1_18/Y in_wai OAI21X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6734 vdd INVX2_22/Y OAI21X1_18/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6735 gnd INVX2_10/Y OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6736 OAI21X1_18/a_2_6# in_wai gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6737 OAI21X1_18/Y INVX2_22/Y OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6738 OAI21X1_16/a_9_54# INVX2_10/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6739 AOI21X1_2/B OAI21X1_28/A OAI21X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6740 vdd INVX2_21/A AOI21X1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6741 gnd INVX2_10/Y OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6742 OAI21X1_16/a_2_6# OAI21X1_28/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6743 AOI21X1_2/B INVX2_21/A OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6744 NOR2X1_4/a_9_54# in_wai vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6745 NOR2X1_4/Y con_loseSig NOR2X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6746 NOR2X1_4/Y in_wai gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6747 gnd con_loseSig NOR2X1_4/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6748 NAND3X1_6/Y in_run vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6749 vdd INVX2_21/Y NAND3X1_6/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6750 NAND3X1_6/Y NOR2X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6751 NAND3X1_6/a_9_6# in_run gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6752 NAND3X1_6/a_14_6# INVX2_21/Y NAND3X1_6/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6753 NAND3X1_6/Y NOR2X1_4/Y NAND3X1_6/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6754 NAND2X1_6/Y con_loseSig vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6755 vdd INVX2_21/Y NAND2X1_6/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6756 NAND2X1_6/a_9_6# con_loseSig gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6757 NAND2X1_6/Y INVX2_21/Y NAND2X1_6/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6758 NAND3X1_5/Y INVX2_8/Y vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6759 vdd INVX2_18/Y NAND3X1_5/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6760 NAND3X1_5/Y INVX2_20/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6761 NAND3X1_5/a_9_6# INVX2_8/Y gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6762 NAND3X1_5/a_14_6# INVX2_18/Y NAND3X1_5/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6763 NAND3X1_5/Y INVX2_20/Y NAND3X1_5/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6764 INVX2_18/Y in_wai vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6765 INVX2_18/Y in_wai gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6766 vdd INVX2_30/A XOR2X1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6767 XOR2X1_25/a_18_54# XOR2X1_25/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6768 OAI21X1_6/B INVX2_30/A XOR2X1_25/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6769 XOR2X1_25/a_35_54# XOR2X1_25/a_2_6# OAI21X1_6/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6770 vdd NOR2X1_3/B XOR2X1_25/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6771 XOR2X1_25/a_13_43# NOR2X1_3/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6772 gnd INVX2_30/A XOR2X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6773 XOR2X1_25/a_18_6# XOR2X1_25/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6774 OAI21X1_6/B XOR2X1_25/a_2_6# XOR2X1_25/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6775 XOR2X1_25/a_35_6# INVX2_30/A OAI21X1_6/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6776 gnd NOR2X1_3/B XOR2X1_25/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6777 XOR2X1_25/a_13_43# NOR2X1_3/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6778 NOR2X1_3/a_9_54# INVX2_30/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6779 NOR2X1_3/Y NOR2X1_3/B NOR2X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6780 NOR2X1_3/Y INVX2_30/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M6781 gnd NOR2X1_3/B NOR2X1_3/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6782 vdd XOR2X1_24/A XOR2X1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6783 XOR2X1_24/a_18_54# XOR2X1_24/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6784 XOR2X1_24/Y XOR2X1_24/A XOR2X1_24/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6785 XOR2X1_24/a_35_54# XOR2X1_24/a_2_6# XOR2X1_24/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6786 vdd NOR2X1_3/Y XOR2X1_24/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6787 XOR2X1_24/a_13_43# NOR2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6788 gnd XOR2X1_24/A XOR2X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6789 XOR2X1_24/a_18_6# XOR2X1_24/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6790 XOR2X1_24/Y XOR2X1_24/a_2_6# XOR2X1_24/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6791 XOR2X1_24/a_35_6# XOR2X1_24/A XOR2X1_24/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6792 gnd NOR2X1_3/Y XOR2X1_24/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6793 XOR2X1_24/a_13_43# NOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6794 vdd XOR2X1_23/A AOI22X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6795 AOI22X1_16/a_2_54# out_MuxData[14] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6796 NOR2X1_3/B out_MuxData[13] AOI22X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6797 AOI22X1_16/a_2_54# XOR2X1_22/A NOR2X1_3/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6798 AOI22X1_16/a_11_6# XOR2X1_23/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6799 NOR2X1_3/B out_MuxData[14] AOI22X1_16/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6800 AOI22X1_16/a_28_6# out_MuxData[13] NOR2X1_3/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6801 gnd XOR2X1_22/A AOI22X1_16/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6802 vdd XOR2X1_23/A XOR2X1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6803 XOR2X1_23/a_18_54# XOR2X1_23/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6804 XOR2X1_22/A XOR2X1_23/A XOR2X1_23/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6805 XOR2X1_23/a_35_54# XOR2X1_23/a_2_6# XOR2X1_22/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6806 vdd out_MuxData[14] XOR2X1_23/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6807 XOR2X1_23/a_13_43# out_MuxData[14] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6808 gnd XOR2X1_23/A XOR2X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6809 XOR2X1_23/a_18_6# XOR2X1_23/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6810 XOR2X1_22/A XOR2X1_23/a_2_6# XOR2X1_23/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6811 XOR2X1_23/a_35_6# XOR2X1_23/A XOR2X1_22/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6812 gnd out_MuxData[14] XOR2X1_23/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6813 XOR2X1_23/a_13_43# out_MuxData[14] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6814 vdd XNOR2X1_3/Y AOI22X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M6815 AOI22X1_15/a_2_54# INVX2_26/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6816 AND2X2_17/A INVX2_25/Y AOI22X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M6817 AOI22X1_15/a_2_54# XNOR2X1_5/Y AND2X2_17/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6818 AOI22X1_15/a_11_6# XNOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6819 AND2X2_17/A INVX2_26/Y AOI22X1_15/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6820 AOI22X1_15/a_28_6# INVX2_25/Y AND2X2_17/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6821 gnd XNOR2X1_5/Y AOI22X1_15/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6822 INVX2_17/Y out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6823 INVX2_17/Y out_MuxData[7] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6824 NAND2X1_5/Y out_MuxData[12] vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6825 vdd out_MuxData[13] NAND2X1_5/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6826 NAND2X1_5/a_9_6# out_MuxData[12] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6827 NAND2X1_5/Y out_MuxData[13] NAND2X1_5/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6828 OAI21X1_14/a_9_54# INVX2_5/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6829 INVX2_27/A XNOR2X1_9/A OAI21X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6830 vdd NAND2X1_5/Y INVX2_27/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6831 gnd INVX2_5/A OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6832 OAI21X1_14/a_2_6# XNOR2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6833 INVX2_27/A NAND2X1_5/Y OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6834 OAI21X1_12/a_9_54# out_MuxData[13] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6835 XNOR2X1_9/A out_MuxData[12] OAI21X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6836 vdd NAND2X1_5/Y XNOR2X1_9/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6837 gnd out_MuxData[13] OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6838 OAI21X1_12/a_2_6# out_MuxData[12] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6839 XNOR2X1_9/A NAND2X1_5/Y OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6840 vdd NOR2X1_8/B XNOR2X1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6841 XNOR2X1_10/a_18_54# XNOR2X1_10/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6842 NAND2X1_4/B XNOR2X1_10/a_2_6# XNOR2X1_10/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6843 XNOR2X1_10/a_35_54# NOR2X1_8/B NAND2X1_4/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6844 vdd NOR2X1_8/A XNOR2X1_10/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6845 XNOR2X1_10/a_12_41# NOR2X1_8/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6846 gnd NOR2X1_8/B XNOR2X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6847 XNOR2X1_10/a_18_6# XNOR2X1_10/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6848 NAND2X1_4/B NOR2X1_8/B XNOR2X1_10/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6849 XNOR2X1_10/a_35_6# XNOR2X1_10/a_2_6# NAND2X1_4/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6850 gnd NOR2X1_8/A XNOR2X1_10/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6851 XNOR2X1_10/a_12_41# NOR2X1_8/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6852 vdd out_MuxData[12] XOR2X1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6853 XOR2X1_18/a_18_54# XOR2X1_18/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6854 AND2X2_8/B out_MuxData[12] XOR2X1_18/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6855 XOR2X1_18/a_35_54# XOR2X1_18/a_2_6# AND2X2_8/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6856 vdd XOR2X1_18/B XOR2X1_18/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6857 XOR2X1_18/a_13_43# XOR2X1_18/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6858 gnd out_MuxData[12] XOR2X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6859 XOR2X1_18/a_18_6# XOR2X1_18/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6860 AND2X2_8/B XOR2X1_18/a_2_6# XOR2X1_18/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6861 XOR2X1_18/a_35_6# out_MuxData[12] AND2X2_8/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6862 gnd XOR2X1_18/B XOR2X1_18/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6863 XOR2X1_18/a_13_43# XOR2X1_18/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6864 OAI21X1_11/a_9_54# NAND2X1_4/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6865 XOR2X1_27/A NAND2X1_4/B OAI21X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6866 vdd NAND3X1_3/Y XOR2X1_27/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6867 gnd NAND2X1_4/A OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6868 OAI21X1_11/a_2_6# NAND2X1_4/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6869 XOR2X1_27/A NAND3X1_3/Y OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6870 NAND3X1_3/Y AND2X2_14/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M6871 vdd NAND2X1_4/Y NAND3X1_3/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6872 NAND3X1_3/Y NAND3X1_3/C vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6873 NAND3X1_3/a_9_6# AND2X2_14/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6874 NAND3X1_3/a_14_6# NAND2X1_4/Y NAND3X1_3/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M6875 NAND3X1_3/Y NAND3X1_3/C NAND3X1_3/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M6876 NAND2X1_4/Y NAND2X1_4/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6877 vdd NAND2X1_4/B NAND2X1_4/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6878 NAND2X1_4/a_9_6# NAND2X1_4/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6879 NAND2X1_4/Y NAND2X1_4/B NAND2X1_4/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6880 OAI21X1_10/a_9_54# NAND2X1_4/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6881 XNOR2X1_8/A NAND2X1_4/B OAI21X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6882 vdd NAND2X1_4/Y XNOR2X1_8/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6883 gnd NAND2X1_4/A OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6884 OAI21X1_10/a_2_6# NAND2X1_4/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6885 XNOR2X1_8/A NAND2X1_4/Y OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6886 vdd XNOR2X1_8/A XNOR2X1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6887 XNOR2X1_8/a_18_54# XNOR2X1_8/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6888 XNOR2X1_8/Y XNOR2X1_8/a_2_6# XNOR2X1_8/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6889 XNOR2X1_8/a_35_54# XNOR2X1_8/A XNOR2X1_8/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6890 vdd AND2X2_14/Y XNOR2X1_8/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6891 XNOR2X1_8/a_12_41# AND2X2_14/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6892 gnd XNOR2X1_8/A XNOR2X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6893 XNOR2X1_8/a_18_6# XNOR2X1_8/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6894 XNOR2X1_8/Y XNOR2X1_8/A XNOR2X1_8/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6895 XNOR2X1_8/a_35_6# XNOR2X1_8/a_2_6# XNOR2X1_8/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6896 gnd AND2X2_14/Y XNOR2X1_8/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6897 XNOR2X1_8/a_12_41# AND2X2_14/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6898 vdd XNOR2X1_7/A XNOR2X1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6899 XNOR2X1_7/a_18_54# XNOR2X1_7/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6900 XNOR2X1_7/Y XNOR2X1_7/a_2_6# XNOR2X1_7/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M6901 XNOR2X1_7/a_35_54# XNOR2X1_7/A XNOR2X1_7/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6902 vdd AND2X2_8/Y XNOR2X1_7/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6903 XNOR2X1_7/a_12_41# AND2X2_8/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6904 gnd XNOR2X1_7/A XNOR2X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6905 XNOR2X1_7/a_18_6# XNOR2X1_7/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6906 XNOR2X1_7/Y XNOR2X1_7/A XNOR2X1_7/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M6907 XNOR2X1_7/a_35_6# XNOR2X1_7/a_2_6# XNOR2X1_7/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6908 gnd AND2X2_8/Y XNOR2X1_7/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6909 XNOR2X1_7/a_12_41# AND2X2_8/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6910 AND2X2_8/a_2_6# AND2X2_8/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6911 vdd AND2X2_8/B AND2X2_8/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6912 AND2X2_8/Y AND2X2_8/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6913 AND2X2_8/a_9_6# AND2X2_8/A AND2X2_8/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6914 gnd AND2X2_8/B AND2X2_8/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6915 AND2X2_8/Y AND2X2_8/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6916 vdd INVX2_41/Y DFFPOSX1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6917 DFFPOSX1_13/a_17_74# INVX2_24/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6918 DFFPOSX1_13/a_22_6# INVX2_41/Y DFFPOSX1_13/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6919 DFFPOSX1_13/a_31_74# DFFPOSX1_13/a_2_6# DFFPOSX1_13/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6920 vdd DFFPOSX1_13/a_34_4# DFFPOSX1_13/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6921 DFFPOSX1_13/a_34_4# DFFPOSX1_13/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6922 DFFPOSX1_13/a_61_74# DFFPOSX1_13/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6923 DFFPOSX1_13/a_66_6# DFFPOSX1_13/a_2_6# DFFPOSX1_13/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6924 DFFPOSX1_13/a_76_84# INVX2_41/Y DFFPOSX1_13/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6925 vdd con_countWriteout[2] DFFPOSX1_13/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6926 gnd INVX2_41/Y DFFPOSX1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6927 con_countWriteout[2] DFFPOSX1_13/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6928 DFFPOSX1_13/a_17_6# INVX2_24/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6929 DFFPOSX1_13/a_22_6# DFFPOSX1_13/a_2_6# DFFPOSX1_13/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6930 DFFPOSX1_13/a_31_6# INVX2_41/Y DFFPOSX1_13/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6931 gnd DFFPOSX1_13/a_34_4# DFFPOSX1_13/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6932 DFFPOSX1_13/a_34_4# DFFPOSX1_13/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6933 DFFPOSX1_13/a_61_6# DFFPOSX1_13/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6934 DFFPOSX1_13/a_66_6# INVX2_41/Y DFFPOSX1_13/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6935 DFFPOSX1_13/a_76_6# DFFPOSX1_13/a_2_6# DFFPOSX1_13/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6936 gnd con_countWriteout[2] DFFPOSX1_13/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6937 con_countWriteout[2] DFFPOSX1_13/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6938 vdd BUFX2_5/Y DFFPOSX1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6939 DFFPOSX1_12/a_17_74# AND2X2_7/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6940 DFFPOSX1_12/a_22_6# BUFX2_5/Y DFFPOSX1_12/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6941 DFFPOSX1_12/a_31_74# DFFPOSX1_12/a_2_6# DFFPOSX1_12/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6942 vdd DFFPOSX1_12/a_34_4# DFFPOSX1_12/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6943 DFFPOSX1_12/a_34_4# DFFPOSX1_12/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6944 DFFPOSX1_12/a_61_74# DFFPOSX1_12/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6945 DFFPOSX1_12/a_66_6# DFFPOSX1_12/a_2_6# DFFPOSX1_12/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6946 DFFPOSX1_12/a_76_84# BUFX2_5/Y DFFPOSX1_12/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6947 vdd AOI22X1_10/C DFFPOSX1_12/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6948 gnd BUFX2_5/Y DFFPOSX1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6949 AOI22X1_10/C DFFPOSX1_12/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6950 DFFPOSX1_12/a_17_6# AND2X2_7/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6951 DFFPOSX1_12/a_22_6# DFFPOSX1_12/a_2_6# DFFPOSX1_12/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6952 DFFPOSX1_12/a_31_6# BUFX2_5/Y DFFPOSX1_12/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6953 gnd DFFPOSX1_12/a_34_4# DFFPOSX1_12/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6954 DFFPOSX1_12/a_34_4# DFFPOSX1_12/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6955 DFFPOSX1_12/a_61_6# DFFPOSX1_12/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6956 DFFPOSX1_12/a_66_6# BUFX2_5/Y DFFPOSX1_12/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6957 DFFPOSX1_12/a_76_6# DFFPOSX1_12/a_2_6# DFFPOSX1_12/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6958 gnd AOI22X1_10/C DFFPOSX1_12/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6959 AOI22X1_10/C DFFPOSX1_12/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6960 AND2X2_7/a_2_6# HAX1_4/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6961 vdd AND2X2_6/B AND2X2_7/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6962 AND2X2_7/Y AND2X2_7/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6963 AND2X2_7/a_9_6# HAX1_4/YS AND2X2_7/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M6964 gnd AND2X2_6/B AND2X2_7/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6965 AND2X2_7/Y AND2X2_7/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6966 OAI21X1_9/a_9_54# con_countWriteout[1] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M6967 OAI21X1_9/Y con_countWriteout[2] OAI21X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M6968 vdd con_countWriteout[4] OAI21X1_9/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6969 gnd con_countWriteout[1] OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M6970 OAI21X1_9/a_2_6# con_countWriteout[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6971 OAI21X1_9/Y con_countWriteout[4] OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6972 INVX2_12/Y INVX2_12/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6973 INVX2_12/Y INVX2_12/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6974 vdd INVX2_41/Y DFFPOSX1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M6975 DFFPOSX1_11/a_17_74# INVX2_12/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6976 DFFPOSX1_11/a_22_6# INVX2_41/Y DFFPOSX1_11/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M6977 DFFPOSX1_11/a_31_74# DFFPOSX1_11/a_2_6# DFFPOSX1_11/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M6978 vdd DFFPOSX1_11/a_34_4# DFFPOSX1_11/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6979 DFFPOSX1_11/a_34_4# DFFPOSX1_11/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6980 DFFPOSX1_11/a_61_74# DFFPOSX1_11/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M6981 DFFPOSX1_11/a_66_6# DFFPOSX1_11/a_2_6# DFFPOSX1_11/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M6982 DFFPOSX1_11/a_76_84# INVX2_41/Y DFFPOSX1_11/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6983 vdd con_countWriteout[1] DFFPOSX1_11/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6984 gnd INVX2_41/Y DFFPOSX1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M6985 con_countWriteout[1] DFFPOSX1_11/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6986 DFFPOSX1_11/a_17_6# INVX2_12/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6987 DFFPOSX1_11/a_22_6# DFFPOSX1_11/a_2_6# DFFPOSX1_11/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6988 DFFPOSX1_11/a_31_6# INVX2_41/Y DFFPOSX1_11/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6989 gnd DFFPOSX1_11/a_34_4# DFFPOSX1_11/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6990 DFFPOSX1_11/a_34_4# DFFPOSX1_11/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M6991 DFFPOSX1_11/a_61_6# DFFPOSX1_11/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6992 DFFPOSX1_11/a_66_6# INVX2_41/Y DFFPOSX1_11/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M6993 DFFPOSX1_11/a_76_6# DFFPOSX1_11/a_2_6# DFFPOSX1_11/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M6994 gnd con_countWriteout[1] DFFPOSX1_11/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6995 con_countWriteout[1] DFFPOSX1_11/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6996 INVX2_11/Y INVX2_11/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6997 INVX2_11/Y INVX2_11/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M6998 INVX2_10/Y INVX2_10/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M6999 INVX2_10/Y INVX2_10/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7000 vdd in_wai AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M7001 AOI21X1_2/a_2_54# AOI21X1_2/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7002 AOI21X1_2/Y OAI21X1_7/Y AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7003 AOI21X1_2/a_12_6# in_wai gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7004 AOI21X1_2/Y AOI21X1_2/B AOI21X1_2/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M7005 gnd OAI21X1_7/Y AOI21X1_2/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7006 vdd BUFX2_5/Y DFFPOSX1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7007 DFFPOSX1_9/a_17_74# AND2X2_6/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7008 DFFPOSX1_9/a_22_6# BUFX2_5/Y DFFPOSX1_9/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7009 DFFPOSX1_9/a_31_74# DFFPOSX1_9/a_2_6# DFFPOSX1_9/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7010 vdd DFFPOSX1_9/a_34_4# DFFPOSX1_9/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7011 DFFPOSX1_9/a_34_4# DFFPOSX1_9/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7012 DFFPOSX1_9/a_61_74# DFFPOSX1_9/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7013 DFFPOSX1_9/a_66_6# DFFPOSX1_9/a_2_6# DFFPOSX1_9/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7014 DFFPOSX1_9/a_76_84# BUFX2_5/Y DFFPOSX1_9/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7015 vdd AOI22X1_9/C DFFPOSX1_9/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7016 gnd BUFX2_5/Y DFFPOSX1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7017 AOI22X1_9/C DFFPOSX1_9/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7018 DFFPOSX1_9/a_17_6# AND2X2_6/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7019 DFFPOSX1_9/a_22_6# DFFPOSX1_9/a_2_6# DFFPOSX1_9/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7020 DFFPOSX1_9/a_31_6# BUFX2_5/Y DFFPOSX1_9/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7021 gnd DFFPOSX1_9/a_34_4# DFFPOSX1_9/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7022 DFFPOSX1_9/a_34_4# DFFPOSX1_9/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7023 DFFPOSX1_9/a_61_6# DFFPOSX1_9/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7024 DFFPOSX1_9/a_66_6# BUFX2_5/Y DFFPOSX1_9/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7025 DFFPOSX1_9/a_76_6# DFFPOSX1_9/a_2_6# DFFPOSX1_9/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7026 gnd AOI22X1_9/C DFFPOSX1_9/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7027 AOI22X1_9/C DFFPOSX1_9/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7028 OAI21X1_7/a_9_54# INVX2_8/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7029 OAI21X1_7/Y NAND2X1_6/Y OAI21X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7030 vdd INVX2_19/A OAI21X1_7/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7031 gnd INVX2_8/Y OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7032 OAI21X1_7/a_2_6# NAND2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7033 OAI21X1_7/Y INVX2_19/A OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7034 INVX2_8/Y in_run vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7035 INVX2_8/Y in_run gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7036 OAI21X1_15/a_9_54# NAND2X1_3/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7037 XOR2X1_24/A OAI21X1_6/B OAI21X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7038 vdd NAND3X1_4/Y XOR2X1_24/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7039 gnd NAND2X1_3/A OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7040 OAI21X1_15/a_2_6# OAI21X1_6/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7041 XOR2X1_24/A NAND3X1_4/Y OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7042 NAND3X1_4/Y AND2X2_9/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M7043 vdd NAND3X1_4/B NAND3X1_4/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7044 NAND3X1_4/Y AND2X2_9/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7045 NAND3X1_4/a_9_6# AND2X2_9/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7046 NAND3X1_4/a_14_6# NAND3X1_4/B NAND3X1_4/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7047 NAND3X1_4/Y AND2X2_9/B NAND3X1_4/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M7048 vdd XOR2X1_22/A XOR2X1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7049 XOR2X1_22/a_18_54# XOR2X1_22/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7050 AND2X2_9/A XOR2X1_22/A XOR2X1_22/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7051 XOR2X1_22/a_35_54# XOR2X1_22/a_2_6# AND2X2_9/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7052 vdd out_MuxData[13] XOR2X1_22/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7053 XOR2X1_22/a_13_43# out_MuxData[13] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7054 gnd XOR2X1_22/A XOR2X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7055 XOR2X1_22/a_18_6# XOR2X1_22/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7056 AND2X2_9/A XOR2X1_22/a_2_6# XOR2X1_22/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7057 XOR2X1_22/a_35_6# XOR2X1_22/A AND2X2_9/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7058 gnd out_MuxData[13] XOR2X1_22/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7059 XOR2X1_22/a_13_43# out_MuxData[13] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7060 AND2X2_9/a_2_6# AND2X2_9/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7061 vdd AND2X2_9/B AND2X2_9/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7062 AND2X2_9/Y AND2X2_9/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7063 AND2X2_9/a_9_6# AND2X2_9/A AND2X2_9/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7064 gnd AND2X2_9/B AND2X2_9/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7065 AND2X2_9/Y AND2X2_9/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7066 vdd AND2X2_9/A XOR2X1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7067 XOR2X1_21/a_18_54# XOR2X1_21/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7068 XOR2X1_21/Y AND2X2_9/A XOR2X1_21/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7069 XOR2X1_21/a_35_54# XOR2X1_21/a_2_6# XOR2X1_21/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7070 vdd AND2X2_9/B XOR2X1_21/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7071 XOR2X1_21/a_13_43# AND2X2_9/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7072 gnd AND2X2_9/A XOR2X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7073 XOR2X1_21/a_18_6# XOR2X1_21/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7074 XOR2X1_21/Y XOR2X1_21/a_2_6# XOR2X1_21/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7075 XOR2X1_21/a_35_6# AND2X2_9/A XOR2X1_21/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7076 gnd AND2X2_9/B XOR2X1_21/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7077 XOR2X1_21/a_13_43# AND2X2_9/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7078 vdd out_MuxData[4] XOR2X1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7079 XOR2X1_20/a_18_54# XOR2X1_20/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7080 AND2X2_5/B out_MuxData[4] XOR2X1_20/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7081 XOR2X1_20/a_35_54# XOR2X1_20/a_2_6# AND2X2_5/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7082 vdd XOR2X1_30/Y XOR2X1_20/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7083 XOR2X1_20/a_13_43# XOR2X1_30/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7084 gnd out_MuxData[4] XOR2X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7085 XOR2X1_20/a_18_6# XOR2X1_20/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7086 AND2X2_5/B XOR2X1_20/a_2_6# XOR2X1_20/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7087 XOR2X1_20/a_35_6# out_MuxData[4] AND2X2_5/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7088 gnd XOR2X1_30/Y XOR2X1_20/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7089 XOR2X1_20/a_13_43# XOR2X1_30/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7090 vdd INVX2_25/Y AOI22X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7091 AOI22X1_14/a_2_54# XOR2X1_21/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7092 NAND3X1_16/B XOR2X1_11/Y AOI22X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7093 AOI22X1_14/a_2_54# INVX2_26/Y NAND3X1_16/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7094 AOI22X1_14/a_11_6# INVX2_25/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7095 NAND3X1_16/B XOR2X1_21/Y AOI22X1_14/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7096 AOI22X1_14/a_28_6# XOR2X1_11/Y NAND3X1_16/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7097 gnd INVX2_26/Y AOI22X1_14/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7098 vdd out_MuxData[6] AOI22X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7099 AOI22X1_13/a_2_54# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7100 NOR2X1_2/A out_MuxData[2] AOI22X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7101 AOI22X1_13/a_2_54# XOR2X1_19/Y NOR2X1_2/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7102 AOI22X1_13/a_11_6# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7103 NOR2X1_2/A out_MuxData[7] AOI22X1_13/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7104 AOI22X1_13/a_28_6# out_MuxData[2] NOR2X1_2/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7105 gnd XOR2X1_19/Y AOI22X1_13/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7106 vdd INVX2_16/Y XOR2X1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7107 XOR2X1_19/a_18_54# XOR2X1_19/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7108 XOR2X1_19/Y INVX2_16/Y XOR2X1_19/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7109 XOR2X1_19/a_35_54# XOR2X1_19/a_2_6# XOR2X1_19/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7110 vdd INVX2_17/Y XOR2X1_19/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7111 XOR2X1_19/a_13_43# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7112 gnd INVX2_16/Y XOR2X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7113 XOR2X1_19/a_18_6# XOR2X1_19/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7114 XOR2X1_19/Y XOR2X1_19/a_2_6# XOR2X1_19/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7115 XOR2X1_19/a_35_6# INVX2_16/Y XOR2X1_19/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7116 gnd INVX2_17/Y XOR2X1_19/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7117 XOR2X1_19/a_13_43# INVX2_17/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7118 INVX2_16/Y out_MuxData[6] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7119 INVX2_16/Y out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7120 OAI21X1_13/a_9_54# XOR2X1_17/B vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7121 INVX2_4/A XNOR2X1_9/A OAI21X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7122 vdd NAND2X1_5/Y INVX2_4/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7123 gnd XOR2X1_17/B OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7124 OAI21X1_13/a_2_6# XNOR2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7125 INVX2_4/A NAND2X1_5/Y OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7126 vdd XNOR2X1_9/A XNOR2X1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7127 XNOR2X1_9/a_18_54# XNOR2X1_9/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7128 XOR2X1_6/A XNOR2X1_9/a_2_6# XNOR2X1_9/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7129 XNOR2X1_9/a_35_54# XNOR2X1_9/A XOR2X1_6/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7130 vdd out_MuxData[8] XNOR2X1_9/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7131 XNOR2X1_9/a_12_41# out_MuxData[8] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7132 gnd XNOR2X1_9/A XNOR2X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7133 XNOR2X1_9/a_18_6# XNOR2X1_9/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7134 XOR2X1_6/A XNOR2X1_9/A XNOR2X1_9/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7135 XNOR2X1_9/a_35_6# XNOR2X1_9/a_2_6# XOR2X1_6/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7136 gnd out_MuxData[8] XNOR2X1_9/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7137 XNOR2X1_9/a_12_41# out_MuxData[8] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7138 vdd INVX2_16/Y XOR2X1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7139 XOR2X1_17/a_18_54# XOR2X1_17/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7140 XOR2X1_18/B INVX2_16/Y XOR2X1_17/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7141 XOR2X1_17/a_35_54# XOR2X1_17/a_2_6# XOR2X1_18/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7142 vdd XOR2X1_17/B XOR2X1_17/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7143 XOR2X1_17/a_13_43# XOR2X1_17/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7144 gnd INVX2_16/Y XOR2X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7145 XOR2X1_17/a_18_6# XOR2X1_17/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7146 XOR2X1_18/B XOR2X1_17/a_2_6# XOR2X1_17/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7147 XOR2X1_17/a_35_6# INVX2_16/Y XOR2X1_18/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7148 gnd XOR2X1_17/B XOR2X1_17/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7149 XOR2X1_17/a_13_43# XOR2X1_17/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7150 vdd out_MuxData[6] AOI22X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7151 AOI22X1_12/a_2_54# out_MuxData[8] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7152 OAI21X1_0/A out_MuxData[12] AOI22X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7153 AOI22X1_12/a_2_54# XOR2X1_18/B OAI21X1_0/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7154 AOI22X1_12/a_11_6# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7155 OAI21X1_0/A out_MuxData[8] AOI22X1_12/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7156 AOI22X1_12/a_28_6# out_MuxData[12] OAI21X1_0/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7157 gnd XOR2X1_18/B AOI22X1_12/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7158 vdd INVX2_28/Y XOR2X1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7159 XOR2X1_16/a_18_54# XOR2X1_16/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7160 XOR2X1_15/B INVX2_28/Y XOR2X1_16/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7161 XOR2X1_16/a_35_54# XOR2X1_16/a_2_6# XOR2X1_15/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7162 vdd INVX2_5/A XOR2X1_16/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7163 XOR2X1_16/a_13_43# INVX2_5/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7164 gnd INVX2_28/Y XOR2X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7165 XOR2X1_16/a_18_6# XOR2X1_16/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7166 XOR2X1_15/B XOR2X1_16/a_2_6# XOR2X1_16/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7167 XOR2X1_16/a_35_6# INVX2_28/Y XOR2X1_15/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7168 gnd INVX2_5/A XOR2X1_16/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7169 XOR2X1_16/a_13_43# INVX2_5/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7170 vdd out_MuxData[10] XOR2X1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7171 XOR2X1_15/a_18_54# XOR2X1_15/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7172 XOR2X1_14/B out_MuxData[10] XOR2X1_15/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7173 XOR2X1_15/a_35_54# XOR2X1_15/a_2_6# XOR2X1_14/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7174 vdd XOR2X1_15/B XOR2X1_15/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7175 XOR2X1_15/a_13_43# XOR2X1_15/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7176 gnd out_MuxData[10] XOR2X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7177 XOR2X1_15/a_18_6# XOR2X1_15/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7178 XOR2X1_14/B XOR2X1_15/a_2_6# XOR2X1_15/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7179 XOR2X1_15/a_35_6# out_MuxData[10] XOR2X1_14/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7180 gnd XOR2X1_15/B XOR2X1_15/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7181 XOR2X1_15/a_13_43# XOR2X1_15/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7182 vdd XNOR2X1_6/B AOI22X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7183 AOI22X1_11/a_2_54# out_MuxData[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7184 NOR2X1_0/B out_MuxData[4] AOI22X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7185 AOI22X1_11/a_2_54# XOR2X1_14/B NOR2X1_0/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7186 AOI22X1_11/a_11_6# XNOR2X1_6/B gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7187 NOR2X1_0/B out_MuxData[7] AOI22X1_11/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7188 AOI22X1_11/a_28_6# out_MuxData[4] NOR2X1_0/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7189 gnd XOR2X1_14/B AOI22X1_11/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7190 vdd out_MuxData[4] XOR2X1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7191 XOR2X1_14/a_18_54# XOR2X1_14/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7192 XNOR2X1_6/B out_MuxData[4] XOR2X1_14/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7193 XOR2X1_14/a_35_54# XOR2X1_14/a_2_6# XNOR2X1_6/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7194 vdd XOR2X1_14/B XOR2X1_14/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7195 XOR2X1_14/a_13_43# XOR2X1_14/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7196 gnd out_MuxData[4] XOR2X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7197 XOR2X1_14/a_18_6# XOR2X1_14/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7198 XNOR2X1_6/B XOR2X1_14/a_2_6# XOR2X1_14/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7199 XOR2X1_14/a_35_6# out_MuxData[4] XNOR2X1_6/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7200 gnd XOR2X1_14/B XOR2X1_14/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7201 XOR2X1_14/a_13_43# XOR2X1_14/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7202 vdd INVX2_17/Y XNOR2X1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7203 XNOR2X1_6/a_18_54# XNOR2X1_6/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7204 AND2X2_8/A XNOR2X1_6/a_2_6# XNOR2X1_6/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7205 XNOR2X1_6/a_35_54# INVX2_17/Y AND2X2_8/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7206 vdd XNOR2X1_6/B XNOR2X1_6/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7207 XNOR2X1_6/a_12_41# XNOR2X1_6/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7208 gnd INVX2_17/Y XNOR2X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7209 XNOR2X1_6/a_18_6# XNOR2X1_6/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7210 AND2X2_8/A INVX2_17/Y XNOR2X1_6/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7211 XNOR2X1_6/a_35_6# XNOR2X1_6/a_2_6# AND2X2_8/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7212 gnd XNOR2X1_6/B XNOR2X1_6/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7213 XNOR2X1_6/a_12_41# XNOR2X1_6/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7214 NAND3X1_2/Y AND2X2_8/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M7215 vdd NAND3X1_2/B NAND3X1_2/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7216 NAND3X1_2/Y AND2X2_8/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7217 NAND3X1_2/a_9_6# AND2X2_8/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7218 NAND3X1_2/a_14_6# NAND3X1_2/B NAND3X1_2/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7219 NAND3X1_2/Y AND2X2_8/B NAND3X1_2/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M7220 vdd AND2X2_8/B XOR2X1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7221 XOR2X1_13/a_18_54# XOR2X1_13/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7222 XOR2X1_13/Y AND2X2_8/B XOR2X1_13/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7223 XOR2X1_13/a_35_54# XOR2X1_13/a_2_6# XOR2X1_13/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7224 vdd AND2X2_8/A XOR2X1_13/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7225 XOR2X1_13/a_13_43# AND2X2_8/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7226 gnd AND2X2_8/B XOR2X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7227 XOR2X1_13/a_18_6# XOR2X1_13/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7228 XOR2X1_13/Y XOR2X1_13/a_2_6# XOR2X1_13/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7229 XOR2X1_13/a_35_6# AND2X2_8/B XOR2X1_13/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7230 gnd AND2X2_8/A XOR2X1_13/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7231 XOR2X1_13/a_13_43# AND2X2_8/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7232 INVX2_15/Y INVX2_15/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7233 INVX2_15/Y INVX2_15/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7234 vdd con_countWriteout[3] AOI22X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7235 AOI22X1_10/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7236 INVX2_15/A INVX2_11/A AOI22X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7237 AOI22X1_10/a_2_54# AOI22X1_10/C INVX2_15/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7238 AOI22X1_10/a_11_6# con_countWriteout[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7239 INVX2_15/A INVX2_11/Y AOI22X1_10/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7240 AOI22X1_10/a_28_6# INVX2_11/A INVX2_15/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7241 gnd AOI22X1_10/C AOI22X1_10/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7242 INVX2_14/Y con_countWriteout[3] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7243 INVX2_14/Y con_countWriteout[3] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7244 vdd con_countWriteout[3] HAX1_4/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M7245 HAX1_4/a_2_74# HAX1_4/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7246 vdd HAX1_4/a_2_74# HAX1_3/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7247 HAX1_4/a_41_74# HAX1_4/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M7248 HAX1_4/a_49_54# HAX1_4/B HAX1_4/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7249 vdd con_countWriteout[3] HAX1_4/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7250 HAX1_4/YS HAX1_4/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7251 HAX1_4/a_9_6# con_countWriteout[3] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7252 HAX1_4/a_2_74# HAX1_4/B HAX1_4/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7253 gnd HAX1_4/a_2_74# HAX1_3/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M7254 HAX1_4/a_38_6# HAX1_4/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M7255 HAX1_4/a_41_74# HAX1_4/B HAX1_4/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7256 HAX1_4/a_38_6# con_countWriteout[3] HAX1_4/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7257 HAX1_4/YS HAX1_4/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7258 INVX2_13/Y con_countWriteout[4] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7259 INVX2_13/Y con_countWriteout[4] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7260 OAI21X1_8/a_9_54# INVX2_14/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7261 OAI21X1_8/Y INVX2_13/Y OAI21X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7262 vdd OAI21X1_9/Y OAI21X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7263 gnd INVX2_14/Y OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7264 OAI21X1_8/a_2_6# INVX2_13/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7265 OAI21X1_8/Y OAI21X1_9/Y OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7266 OAI22X1_0/a_9_54# con_countWriteout[5] vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7267 INVX2_10/A OR2X1_1/Y OAI22X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=480 pd=104 as=0 ps=0
M7268 OAI22X1_0/a_28_54# OAI21X1_8/Y INVX2_10/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7269 vdd OR2X1_1/Y OAI22X1_0/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7270 gnd con_countWriteout[5] OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=320 ps=152
M7271 OAI22X1_0/a_2_6# OR2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7272 INVX2_10/A OAI21X1_8/Y OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7273 OAI22X1_0/a_2_6# OR2X1_1/Y INVX2_10/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7274 OR2X1_1/a_9_54# con_countWriteout[6] OR2X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M7275 vdd OR2X1_1/B OR2X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7276 OR2X1_1/Y OR2X1_1/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7277 OR2X1_1/a_2_54# con_countWriteout[6] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M7278 gnd OR2X1_1/B OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7279 OR2X1_1/Y OR2X1_1/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7280 vdd INVX2_41/Y DFFPOSX1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7281 DFFPOSX1_10/a_17_74# INVX2_9/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7282 DFFPOSX1_10/a_22_6# INVX2_41/Y DFFPOSX1_10/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7283 DFFPOSX1_10/a_31_74# DFFPOSX1_10/a_2_6# DFFPOSX1_10/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7284 vdd DFFPOSX1_10/a_34_4# DFFPOSX1_10/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7285 DFFPOSX1_10/a_34_4# DFFPOSX1_10/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7286 DFFPOSX1_10/a_61_74# DFFPOSX1_10/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7287 DFFPOSX1_10/a_66_6# DFFPOSX1_10/a_2_6# DFFPOSX1_10/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7288 DFFPOSX1_10/a_76_84# INVX2_41/Y DFFPOSX1_10/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7289 vdd con_countWriteout[6] DFFPOSX1_10/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7290 gnd INVX2_41/Y DFFPOSX1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7291 con_countWriteout[6] DFFPOSX1_10/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7292 DFFPOSX1_10/a_17_6# INVX2_9/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7293 DFFPOSX1_10/a_22_6# DFFPOSX1_10/a_2_6# DFFPOSX1_10/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7294 DFFPOSX1_10/a_31_6# INVX2_41/Y DFFPOSX1_10/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7295 gnd DFFPOSX1_10/a_34_4# DFFPOSX1_10/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7296 DFFPOSX1_10/a_34_4# DFFPOSX1_10/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7297 DFFPOSX1_10/a_61_6# DFFPOSX1_10/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7298 DFFPOSX1_10/a_66_6# INVX2_41/Y DFFPOSX1_10/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7299 DFFPOSX1_10/a_76_6# DFFPOSX1_10/a_2_6# DFFPOSX1_10/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7300 gnd con_countWriteout[6] DFFPOSX1_10/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7301 con_countWriteout[6] DFFPOSX1_10/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7302 INVX2_9/Y INVX2_9/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7303 INVX2_9/Y INVX2_9/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7304 vdd HAX1_0/YC XOR2X1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7305 XOR2X1_12/a_18_54# XOR2X1_12/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7306 AND2X2_6/A HAX1_0/YC XOR2X1_12/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7307 XOR2X1_12/a_35_54# XOR2X1_12/a_2_6# AND2X2_6/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7308 vdd con_countWriteout[8] XOR2X1_12/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7309 XOR2X1_12/a_13_43# con_countWriteout[8] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7310 gnd HAX1_0/YC XOR2X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7311 XOR2X1_12/a_18_6# XOR2X1_12/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7312 AND2X2_6/A XOR2X1_12/a_2_6# XOR2X1_12/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7313 XOR2X1_12/a_35_6# HAX1_0/YC AND2X2_6/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7314 gnd con_countWriteout[8] XOR2X1_12/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7315 XOR2X1_12/a_13_43# con_countWriteout[8] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7316 AND2X2_6/a_2_6# AND2X2_6/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7317 vdd AND2X2_6/B AND2X2_6/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7318 AND2X2_6/Y AND2X2_6/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7319 AND2X2_6/a_9_6# AND2X2_6/A AND2X2_6/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7320 gnd AND2X2_6/B AND2X2_6/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7321 AND2X2_6/Y AND2X2_6/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7322 vdd con_countWriteout[8] AOI22X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7323 AOI22X1_9/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7324 INVX2_7/A INVX2_11/A AOI22X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7325 AOI22X1_9/a_2_54# AOI22X1_9/C INVX2_7/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7326 AOI22X1_9/a_11_6# con_countWriteout[8] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7327 INVX2_7/A INVX2_11/Y AOI22X1_9/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7328 AOI22X1_9/a_28_6# INVX2_11/A INVX2_7/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7329 gnd AOI22X1_9/C AOI22X1_9/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7330 INVX2_7/Y INVX2_7/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7331 INVX2_7/Y INVX2_7/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7332 vdd INVX2_41/Y DFFPOSX1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7333 DFFPOSX1_8/a_17_74# INVX2_7/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7334 DFFPOSX1_8/a_22_6# INVX2_41/Y DFFPOSX1_8/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7335 DFFPOSX1_8/a_31_74# DFFPOSX1_8/a_2_6# DFFPOSX1_8/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7336 vdd DFFPOSX1_8/a_34_4# DFFPOSX1_8/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7337 DFFPOSX1_8/a_34_4# DFFPOSX1_8/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7338 DFFPOSX1_8/a_61_74# DFFPOSX1_8/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7339 DFFPOSX1_8/a_66_6# DFFPOSX1_8/a_2_6# DFFPOSX1_8/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7340 DFFPOSX1_8/a_76_84# INVX2_41/Y DFFPOSX1_8/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7341 vdd con_countWriteout[8] DFFPOSX1_8/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7342 gnd INVX2_41/Y DFFPOSX1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7343 con_countWriteout[8] DFFPOSX1_8/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7344 DFFPOSX1_8/a_17_6# INVX2_7/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7345 DFFPOSX1_8/a_22_6# DFFPOSX1_8/a_2_6# DFFPOSX1_8/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7346 DFFPOSX1_8/a_31_6# INVX2_41/Y DFFPOSX1_8/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7347 gnd DFFPOSX1_8/a_34_4# DFFPOSX1_8/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7348 DFFPOSX1_8/a_34_4# DFFPOSX1_8/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7349 DFFPOSX1_8/a_61_6# DFFPOSX1_8/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7350 DFFPOSX1_8/a_66_6# INVX2_41/Y DFFPOSX1_8/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7351 DFFPOSX1_8/a_76_6# DFFPOSX1_8/a_2_6# DFFPOSX1_8/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7352 gnd con_countWriteout[8] DFFPOSX1_8/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7353 con_countWriteout[8] DFFPOSX1_8/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7354 OAI21X1_6/a_9_54# NAND2X1_3/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7355 XNOR2X1_5/A OAI21X1_6/B OAI21X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7356 vdd NAND3X1_4/B XNOR2X1_5/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7357 gnd NAND2X1_3/A OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7358 OAI21X1_6/a_2_6# OAI21X1_6/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7359 XNOR2X1_5/A NAND3X1_4/B OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7360 vdd XNOR2X1_5/A XNOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7361 XNOR2X1_5/a_18_54# XNOR2X1_5/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7362 XNOR2X1_5/Y XNOR2X1_5/a_2_6# XNOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7363 XNOR2X1_5/a_35_54# XNOR2X1_5/A XNOR2X1_5/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7364 vdd AND2X2_9/Y XNOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7365 XNOR2X1_5/a_12_41# AND2X2_9/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7366 gnd XNOR2X1_5/A XNOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7367 XNOR2X1_5/a_18_6# XNOR2X1_5/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7368 XNOR2X1_5/Y XNOR2X1_5/A XNOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7369 XNOR2X1_5/a_35_6# XNOR2X1_5/a_2_6# XNOR2X1_5/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7370 gnd AND2X2_9/Y XNOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7371 XNOR2X1_5/a_12_41# AND2X2_9/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7372 vdd INVX2_16/Y XNOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7373 XNOR2X1_4/a_18_54# XNOR2X1_4/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7374 AND2X2_9/B XNOR2X1_4/a_2_6# XNOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7375 XNOR2X1_4/a_35_54# INVX2_16/Y AND2X2_9/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7376 vdd XOR2X1_8/Y XNOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7377 XNOR2X1_4/a_12_41# XOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7378 gnd INVX2_16/Y XNOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7379 XNOR2X1_4/a_18_6# XNOR2X1_4/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7380 AND2X2_9/B INVX2_16/Y XNOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7381 XNOR2X1_4/a_35_6# XNOR2X1_4/a_2_6# AND2X2_9/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7382 gnd XOR2X1_8/Y XNOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7383 XNOR2X1_4/a_12_41# XOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7384 vdd OAI21X1_5/Y XNOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7385 XNOR2X1_3/a_18_54# XNOR2X1_3/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7386 XNOR2X1_3/Y XNOR2X1_3/a_2_6# XNOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7387 XNOR2X1_3/a_35_54# OAI21X1_5/Y XNOR2X1_3/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7388 vdd AND2X2_5/Y XNOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7389 XNOR2X1_3/a_12_41# AND2X2_5/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7390 gnd OAI21X1_5/Y XNOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7391 XNOR2X1_3/a_18_6# XNOR2X1_3/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7392 XNOR2X1_3/Y OAI21X1_5/Y XNOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7393 XNOR2X1_3/a_35_6# XNOR2X1_3/a_2_6# XNOR2X1_3/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7394 gnd AND2X2_5/Y XNOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7395 XNOR2X1_3/a_12_41# AND2X2_5/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7396 AND2X2_5/a_2_6# AND2X2_5/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7397 vdd AND2X2_5/B AND2X2_5/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7398 AND2X2_5/Y AND2X2_5/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7399 AND2X2_5/a_9_6# AND2X2_5/A AND2X2_5/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7400 gnd AND2X2_5/B AND2X2_5/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7401 AND2X2_5/Y AND2X2_5/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7402 NAND3X1_1/Y AND2X2_5/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M7403 vdd NAND3X1_1/B NAND3X1_1/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7404 NAND3X1_1/Y AND2X2_5/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7405 NAND3X1_1/a_9_6# AND2X2_5/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7406 NAND3X1_1/a_14_6# NAND3X1_1/B NAND3X1_1/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7407 NAND3X1_1/Y AND2X2_5/B NAND3X1_1/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M7408 vdd AND2X2_5/B XOR2X1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7409 XOR2X1_11/a_18_54# XOR2X1_11/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7410 XOR2X1_11/Y AND2X2_5/B XOR2X1_11/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7411 XOR2X1_11/a_35_54# XOR2X1_11/a_2_6# XOR2X1_11/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7412 vdd AND2X2_5/A XOR2X1_11/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7413 XOR2X1_11/a_13_43# AND2X2_5/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7414 gnd AND2X2_5/B XOR2X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7415 XOR2X1_11/a_18_6# XOR2X1_11/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7416 XOR2X1_11/Y XOR2X1_11/a_2_6# XOR2X1_11/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7417 XOR2X1_11/a_35_6# AND2X2_5/B XOR2X1_11/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7418 gnd AND2X2_5/A XOR2X1_11/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7419 XOR2X1_11/a_13_43# AND2X2_5/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7420 vdd out_MuxData[2] XOR2X1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7421 XOR2X1_10/a_18_54# XOR2X1_10/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7422 XOR2X1_9/B out_MuxData[2] XOR2X1_10/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7423 XOR2X1_10/a_35_54# XOR2X1_10/a_2_6# XOR2X1_9/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7424 vdd XOR2X1_19/Y XOR2X1_10/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7425 XOR2X1_10/a_13_43# XOR2X1_19/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7426 gnd out_MuxData[2] XOR2X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7427 XOR2X1_10/a_18_6# XOR2X1_10/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7428 XOR2X1_9/B XOR2X1_10/a_2_6# XOR2X1_10/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7429 XOR2X1_10/a_35_6# out_MuxData[2] XOR2X1_9/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7430 gnd XOR2X1_19/Y XOR2X1_10/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7431 XOR2X1_10/a_13_43# XOR2X1_19/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7432 vdd out_MuxData[12] XOR2X1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7433 XOR2X1_9/a_18_54# XOR2X1_9/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7434 XOR2X1_9/Y out_MuxData[12] XOR2X1_9/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7435 XOR2X1_9/a_35_54# XOR2X1_9/a_2_6# XOR2X1_9/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7436 vdd XOR2X1_9/B XOR2X1_9/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7437 XOR2X1_9/a_13_43# XOR2X1_9/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7438 gnd out_MuxData[12] XOR2X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7439 XOR2X1_9/a_18_6# XOR2X1_9/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7440 XOR2X1_9/Y XOR2X1_9/a_2_6# XOR2X1_9/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7441 XOR2X1_9/a_35_6# out_MuxData[12] XOR2X1_9/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7442 gnd XOR2X1_9/B XOR2X1_9/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7443 XOR2X1_9/a_13_43# XOR2X1_9/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7444 vdd XOR2X1_9/Y AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7445 AOI22X1_7/a_2_54# out_MuxData[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7446 NOR2X1_2/B out_MuxData[12] AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7447 AOI22X1_7/a_2_54# XOR2X1_9/B NOR2X1_2/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7448 AOI22X1_7/a_11_6# XOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7449 NOR2X1_2/B out_MuxData[15] AOI22X1_7/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7450 AOI22X1_7/a_28_6# out_MuxData[12] NOR2X1_2/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7451 gnd XOR2X1_9/B AOI22X1_7/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7452 out_MuxData[15] INVX2_5/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7453 out_MuxData[15] INVX2_5/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7454 vdd XOR2X1_6/A XOR2X1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7455 XOR2X1_6/a_18_54# XOR2X1_6/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7456 XOR2X1_5/A XOR2X1_6/A XOR2X1_6/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7457 XOR2X1_6/a_35_54# XOR2X1_6/a_2_6# XOR2X1_5/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7458 vdd out_MuxData[6] XOR2X1_6/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7459 XOR2X1_6/a_13_43# out_MuxData[6] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7460 gnd XOR2X1_6/A XOR2X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7461 XOR2X1_6/a_18_6# XOR2X1_6/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7462 XOR2X1_5/A XOR2X1_6/a_2_6# XOR2X1_6/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7463 XOR2X1_6/a_35_6# XOR2X1_6/A XOR2X1_5/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7464 gnd out_MuxData[6] XOR2X1_6/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7465 XOR2X1_6/a_13_43# out_MuxData[6] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7466 vdd XOR2X1_6/A AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7467 AOI22X1_6/a_2_54# out_MuxData[6] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7468 XOR2X1_3/B out_MuxData[5] AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7469 AOI22X1_6/a_2_54# XOR2X1_5/A XOR2X1_3/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7470 AOI22X1_6/a_11_6# XOR2X1_6/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7471 XOR2X1_3/B out_MuxData[6] AOI22X1_6/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7472 AOI22X1_6/a_28_6# out_MuxData[5] XOR2X1_3/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7473 gnd XOR2X1_5/A AOI22X1_6/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7474 vdd XOR2X1_5/A XOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7475 XOR2X1_5/a_18_54# XOR2X1_5/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7476 AND2X2_4/A XOR2X1_5/A XOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7477 XOR2X1_5/a_35_54# XOR2X1_5/a_2_6# AND2X2_4/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7478 vdd out_MuxData[5] XOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7479 XOR2X1_5/a_13_43# out_MuxData[5] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7480 gnd XOR2X1_5/A XOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7481 XOR2X1_5/a_18_6# XOR2X1_5/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7482 AND2X2_4/A XOR2X1_5/a_2_6# XOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7483 XOR2X1_5/a_35_6# XOR2X1_5/A AND2X2_4/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7484 gnd out_MuxData[5] XOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7485 XOR2X1_5/a_13_43# out_MuxData[5] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7486 vdd out_MuxData[4] XOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7487 XOR2X1_4/a_18_54# XOR2X1_4/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7488 XOR2X1_4/Y out_MuxData[4] XOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7489 XOR2X1_4/a_35_54# XOR2X1_4/a_2_6# XOR2X1_4/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7490 vdd out_MuxData[10] XOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7491 XOR2X1_4/a_13_43# out_MuxData[10] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7492 gnd out_MuxData[4] XOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7493 XOR2X1_4/a_18_6# XOR2X1_4/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7494 XOR2X1_4/Y XOR2X1_4/a_2_6# XOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7495 XOR2X1_4/a_35_6# out_MuxData[4] XOR2X1_4/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7496 gnd out_MuxData[10] XOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7497 XOR2X1_4/a_13_43# out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7498 vdd out_MuxData[10] AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7499 AOI22X1_5/a_2_54# out_MuxData[4] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7500 OAI21X1_2/A out_MuxData[14] AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7501 AOI22X1_5/a_2_54# XOR2X1_4/Y OAI21X1_2/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7502 AOI22X1_5/a_11_6# out_MuxData[10] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7503 OAI21X1_2/A out_MuxData[4] AOI22X1_5/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7504 AOI22X1_5/a_28_6# out_MuxData[14] OAI21X1_2/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7505 gnd XOR2X1_4/Y AOI22X1_5/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7506 vdd out_MuxData[14] AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7507 AOI22X1_4/a_2_54# out_MuxData[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7508 NOR2X1_0/A out_MuxData[10] AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7509 AOI22X1_4/a_2_54# XOR2X1_15/B NOR2X1_0/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7510 AOI22X1_4/a_11_6# out_MuxData[14] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7511 NOR2X1_0/A out_MuxData[15] AOI22X1_4/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7512 AOI22X1_4/a_28_6# out_MuxData[10] NOR2X1_0/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7513 gnd XOR2X1_15/B AOI22X1_4/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7514 vdd INVX2_28/Y XNOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7515 XNOR2X1_1/a_18_54# XNOR2X1_1/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7516 XOR2X1_1/B XNOR2X1_1/a_2_6# XNOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7517 XNOR2X1_1/a_35_54# INVX2_28/Y XOR2X1_1/B vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7518 vdd XOR2X1_4/Y XNOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7519 XNOR2X1_1/a_12_41# XOR2X1_4/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7520 gnd INVX2_28/Y XNOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7521 XNOR2X1_1/a_18_6# XNOR2X1_1/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7522 XOR2X1_1/B INVX2_28/Y XNOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7523 XNOR2X1_1/a_35_6# XNOR2X1_1/a_2_6# XOR2X1_1/B Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7524 gnd XOR2X1_4/Y XNOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7525 XNOR2X1_1/a_12_41# XOR2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7526 vdd AND2X2_4/A XOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7527 XOR2X1_1/a_18_54# XOR2X1_1/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7528 XOR2X1_1/Y AND2X2_4/A XOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7529 XOR2X1_1/a_35_54# XOR2X1_1/a_2_6# XOR2X1_1/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7530 vdd XOR2X1_1/B XOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7531 XOR2X1_1/a_13_43# XOR2X1_1/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7532 gnd AND2X2_4/A XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7533 XOR2X1_1/a_18_6# XOR2X1_1/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7534 XOR2X1_1/Y XOR2X1_1/a_2_6# XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7535 XOR2X1_1/a_35_6# AND2X2_4/A XOR2X1_1/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7536 gnd XOR2X1_1/B XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7537 XOR2X1_1/a_13_43# XOR2X1_1/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7538 NOR2X1_0/a_9_54# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7539 XOR2X1_0/B NOR2X1_0/B NOR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7540 XOR2X1_0/B NOR2X1_0/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M7541 gnd NOR2X1_0/B XOR2X1_0/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7542 vdd NOR2X1_0/A AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M7543 AOI21X1_0/a_2_54# NOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7544 INVX2_3/A XOR2X1_0/B AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7545 AOI21X1_0/a_12_6# NOR2X1_0/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7546 INVX2_3/A NOR2X1_0/B AOI21X1_0/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M7547 gnd XOR2X1_0/B INVX2_3/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7548 NAND3X1_2/B OAI21X1_0/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7549 vdd INVX2_3/Y NAND3X1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7550 NAND2X1_0/a_9_6# OAI21X1_0/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7551 NAND3X1_2/B INVX2_3/Y NAND2X1_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7552 OAI21X1_1/a_9_54# OAI21X1_0/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7553 XNOR2X1_7/A INVX2_3/Y OAI21X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7554 vdd NAND3X1_2/B XNOR2X1_7/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7555 gnd OAI21X1_0/A OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7556 OAI21X1_1/a_2_6# INVX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7557 XNOR2X1_7/A NAND3X1_2/B OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7558 vdd INVX2_41/Y DFFPOSX1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7559 DFFPOSX1_7/a_17_74# INVX2_15/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7560 DFFPOSX1_7/a_22_6# INVX2_41/Y DFFPOSX1_7/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7561 DFFPOSX1_7/a_31_74# DFFPOSX1_7/a_2_6# DFFPOSX1_7/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7562 vdd DFFPOSX1_7/a_34_4# DFFPOSX1_7/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7563 DFFPOSX1_7/a_34_4# DFFPOSX1_7/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7564 DFFPOSX1_7/a_61_74# DFFPOSX1_7/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7565 DFFPOSX1_7/a_66_6# DFFPOSX1_7/a_2_6# DFFPOSX1_7/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7566 DFFPOSX1_7/a_76_84# INVX2_41/Y DFFPOSX1_7/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7567 vdd con_countWriteout[3] DFFPOSX1_7/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7568 gnd INVX2_41/Y DFFPOSX1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7569 con_countWriteout[3] DFFPOSX1_7/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7570 DFFPOSX1_7/a_17_6# INVX2_15/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7571 DFFPOSX1_7/a_22_6# DFFPOSX1_7/a_2_6# DFFPOSX1_7/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7572 DFFPOSX1_7/a_31_6# INVX2_41/Y DFFPOSX1_7/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7573 gnd DFFPOSX1_7/a_34_4# DFFPOSX1_7/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7574 DFFPOSX1_7/a_34_4# DFFPOSX1_7/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7575 DFFPOSX1_7/a_61_6# DFFPOSX1_7/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7576 DFFPOSX1_7/a_66_6# INVX2_41/Y DFFPOSX1_7/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7577 DFFPOSX1_7/a_76_6# DFFPOSX1_7/a_2_6# DFFPOSX1_7/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7578 gnd con_countWriteout[3] DFFPOSX1_7/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7579 con_countWriteout[3] DFFPOSX1_7/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7580 INVX2_2/Y INVX2_2/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7581 INVX2_2/Y INVX2_2/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7582 vdd con_countWriteout[4] AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7583 AOI22X1_3/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7584 INVX2_2/A INVX2_11/A AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7585 AOI22X1_3/a_2_54# AOI22X1_3/C INVX2_2/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7586 AOI22X1_3/a_11_6# con_countWriteout[4] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7587 INVX2_2/A INVX2_11/Y AOI22X1_3/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7588 AOI22X1_3/a_28_6# INVX2_11/A INVX2_2/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7589 gnd AOI22X1_3/C AOI22X1_3/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7590 vdd con_countWriteout[4] HAX1_3/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M7591 HAX1_3/a_2_74# HAX1_3/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7592 vdd HAX1_3/a_2_74# HAX1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7593 HAX1_3/a_41_74# HAX1_3/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M7594 HAX1_3/a_49_54# HAX1_3/B HAX1_3/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7595 vdd con_countWriteout[4] HAX1_3/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7596 HAX1_3/YS HAX1_3/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7597 HAX1_3/a_9_6# con_countWriteout[4] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7598 HAX1_3/a_2_74# HAX1_3/B HAX1_3/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7599 gnd HAX1_3/a_2_74# HAX1_2/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M7600 HAX1_3/a_38_6# HAX1_3/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M7601 HAX1_3/a_41_74# HAX1_3/B HAX1_3/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7602 HAX1_3/a_38_6# con_countWriteout[4] HAX1_3/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7603 HAX1_3/YS HAX1_3/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7604 vdd con_countWriteout[5] AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7605 AOI22X1_2/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7606 INVX2_0/A INVX2_11/A AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7607 AOI22X1_2/a_2_54# AOI22X1_2/C INVX2_0/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7608 AOI22X1_2/a_11_6# con_countWriteout[5] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7609 INVX2_0/A INVX2_11/Y AOI22X1_2/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7610 AOI22X1_2/a_28_6# INVX2_11/A INVX2_0/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7611 gnd AOI22X1_2/C AOI22X1_2/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7612 vdd BUFX2_5/Y DFFPOSX1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7613 DFFPOSX1_4/a_17_74# AND2X2_2/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7614 DFFPOSX1_4/a_22_6# BUFX2_5/Y DFFPOSX1_4/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7615 DFFPOSX1_4/a_31_74# DFFPOSX1_4/a_2_6# DFFPOSX1_4/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7616 vdd DFFPOSX1_4/a_34_4# DFFPOSX1_4/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7617 DFFPOSX1_4/a_34_4# DFFPOSX1_4/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7618 DFFPOSX1_4/a_61_74# DFFPOSX1_4/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7619 DFFPOSX1_4/a_66_6# DFFPOSX1_4/a_2_6# DFFPOSX1_4/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7620 DFFPOSX1_4/a_76_84# BUFX2_5/Y DFFPOSX1_4/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7621 vdd AOI22X1_2/C DFFPOSX1_4/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7622 gnd BUFX2_5/Y DFFPOSX1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7623 AOI22X1_2/C DFFPOSX1_4/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7624 DFFPOSX1_4/a_17_6# AND2X2_2/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7625 DFFPOSX1_4/a_22_6# DFFPOSX1_4/a_2_6# DFFPOSX1_4/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7626 DFFPOSX1_4/a_31_6# BUFX2_5/Y DFFPOSX1_4/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7627 gnd DFFPOSX1_4/a_34_4# DFFPOSX1_4/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7628 DFFPOSX1_4/a_34_4# DFFPOSX1_4/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7629 DFFPOSX1_4/a_61_6# DFFPOSX1_4/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7630 DFFPOSX1_4/a_66_6# BUFX2_5/Y DFFPOSX1_4/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7631 DFFPOSX1_4/a_76_6# DFFPOSX1_4/a_2_6# DFFPOSX1_4/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7632 gnd AOI22X1_2/C DFFPOSX1_4/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7633 AOI22X1_2/C DFFPOSX1_4/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7634 vdd con_countWriteout[5] HAX1_2/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M7635 HAX1_2/a_2_74# HAX1_2/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7636 vdd HAX1_2/a_2_74# HAX1_1/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7637 HAX1_2/a_41_74# HAX1_2/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M7638 HAX1_2/a_49_54# HAX1_2/B HAX1_2/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7639 vdd con_countWriteout[5] HAX1_2/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7640 HAX1_2/YS HAX1_2/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7641 HAX1_2/a_9_6# con_countWriteout[5] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7642 HAX1_2/a_2_74# HAX1_2/B HAX1_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7643 gnd HAX1_2/a_2_74# HAX1_1/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M7644 HAX1_2/a_38_6# HAX1_2/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M7645 HAX1_2/a_41_74# HAX1_2/B HAX1_2/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7646 HAX1_2/a_38_6# con_countWriteout[5] HAX1_2/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7647 HAX1_2/YS HAX1_2/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7648 vdd con_countWriteout[6] HAX1_1/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M7649 HAX1_1/a_2_74# HAX1_1/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7650 vdd HAX1_1/a_2_74# HAX1_0/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7651 HAX1_1/a_41_74# HAX1_1/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M7652 HAX1_1/a_49_54# HAX1_1/B HAX1_1/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7653 vdd con_countWriteout[6] HAX1_1/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7654 HAX1_1/YS HAX1_1/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7655 HAX1_1/a_9_6# con_countWriteout[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7656 HAX1_1/a_2_74# HAX1_1/B HAX1_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7657 gnd HAX1_1/a_2_74# HAX1_0/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M7658 HAX1_1/a_38_6# HAX1_1/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M7659 HAX1_1/a_41_74# HAX1_1/B HAX1_1/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7660 HAX1_1/a_38_6# con_countWriteout[6] HAX1_1/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7661 HAX1_1/YS HAX1_1/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7662 vdd con_countWriteout[6] AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7663 AOI22X1_1/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7664 INVX2_9/A INVX2_11/A AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7665 AOI22X1_1/a_2_54# AOI22X1_1/C INVX2_9/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7666 AOI22X1_1/a_11_6# con_countWriteout[6] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7667 INVX2_9/A INVX2_11/Y AOI22X1_1/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7668 AOI22X1_1/a_28_6# INVX2_11/A INVX2_9/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7669 gnd AOI22X1_1/C AOI22X1_1/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7670 OR2X1_0/a_9_54# con_countWriteout[8] OR2X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M7671 vdd con_countWriteout[7] OR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7672 OR2X1_1/B OR2X1_0/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7673 OR2X1_0/a_2_54# con_countWriteout[8] gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M7674 gnd con_countWriteout[7] OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7675 OR2X1_1/B OR2X1_0/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7676 vdd con_countWriteout[7] HAX1_0/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M7677 HAX1_0/a_2_74# HAX1_0/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7678 vdd HAX1_0/a_2_74# HAX1_0/YC vdd pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7679 HAX1_0/a_41_74# HAX1_0/a_2_74# vdd vdd pfet w=20 l=2
+  ad=220 pd=92 as=0 ps=0
M7680 HAX1_0/a_49_54# HAX1_0/B HAX1_0/a_41_74# vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7681 vdd con_countWriteout[7] HAX1_0/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7682 HAX1_0/YS HAX1_0/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7683 HAX1_0/a_9_6# con_countWriteout[7] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7684 HAX1_0/a_2_74# HAX1_0/B HAX1_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7685 gnd HAX1_0/a_2_74# HAX1_0/YC Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M7686 HAX1_0/a_38_6# HAX1_0/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=216 pd=102 as=0 ps=0
M7687 HAX1_0/a_41_74# HAX1_0/B HAX1_0/a_38_6# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7688 HAX1_0/a_38_6# con_countWriteout[7] HAX1_0/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7689 HAX1_0/YS HAX1_0/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7690 vdd con_countWriteout[7] AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7691 AOI22X1_0/a_2_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7692 INVX2_1/A INVX2_11/A AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7693 AOI22X1_0/a_2_54# AOI22X1_0/C INVX2_1/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7694 AOI22X1_0/a_11_6# con_countWriteout[7] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7695 INVX2_1/A INVX2_11/Y AOI22X1_0/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7696 AOI22X1_0/a_28_6# INVX2_11/A INVX2_1/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7697 gnd AOI22X1_0/C AOI22X1_0/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7698 INVX2_1/Y INVX2_1/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7699 INVX2_1/Y INVX2_1/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7700 NAND3X1_4/B NAND2X1_3/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7701 vdd OAI21X1_6/B NAND3X1_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7702 NAND2X1_3/a_9_6# NAND2X1_3/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7703 NAND3X1_4/B OAI21X1_6/B NAND2X1_3/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7704 vdd out_MuxData[2] AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M7705 AOI22X1_8/a_2_54# out_MuxData[12] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7706 NAND2X1_3/A out_MuxData[6] AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M7707 AOI22X1_8/a_2_54# XOR2X1_8/Y NAND2X1_3/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7708 AOI22X1_8/a_11_6# out_MuxData[2] gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7709 NAND2X1_3/A out_MuxData[12] AOI22X1_8/a_11_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7710 AOI22X1_8/a_28_6# out_MuxData[6] NAND2X1_3/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7711 gnd XOR2X1_8/Y AOI22X1_8/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7712 vdd out_MuxData[12] XOR2X1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7713 XOR2X1_8/a_18_54# XOR2X1_8/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7714 XOR2X1_8/Y out_MuxData[12] XOR2X1_8/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7715 XOR2X1_8/a_35_54# XOR2X1_8/a_2_6# XOR2X1_8/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7716 vdd out_MuxData[2] XOR2X1_8/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7717 XOR2X1_8/a_13_43# out_MuxData[2] vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7718 gnd out_MuxData[12] XOR2X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7719 XOR2X1_8/a_18_6# XOR2X1_8/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7720 XOR2X1_8/Y XOR2X1_8/a_2_6# XOR2X1_8/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7721 XOR2X1_8/a_35_6# out_MuxData[12] XOR2X1_8/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7722 gnd out_MuxData[2] XOR2X1_8/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7723 XOR2X1_8/a_13_43# out_MuxData[2] gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7724 OAI21X1_5/a_9_54# OAI21X1_4/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7725 OAI21X1_5/Y INVX2_6/Y OAI21X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7726 vdd NAND3X1_1/B OAI21X1_5/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7727 gnd OAI21X1_4/A OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7728 OAI21X1_5/a_2_6# INVX2_6/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7729 OAI21X1_5/Y NAND3X1_1/B OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7730 NAND3X1_1/B OAI21X1_4/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7731 vdd INVX2_6/Y NAND3X1_1/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7732 NAND2X1_2/a_9_6# OAI21X1_4/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7733 NAND3X1_1/B INVX2_6/Y NAND2X1_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7734 OAI21X1_4/a_9_54# OAI21X1_4/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7735 XOR2X1_7/A INVX2_6/Y OAI21X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7736 vdd NAND3X1_1/Y XOR2X1_7/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7737 gnd OAI21X1_4/A OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7738 OAI21X1_4/a_2_6# INVX2_6/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7739 XOR2X1_7/A NAND3X1_1/Y OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7740 INVX2_6/Y INVX2_6/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7741 INVX2_6/Y INVX2_6/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7742 vdd XOR2X1_7/A XOR2X1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7743 XOR2X1_7/a_18_54# XOR2X1_7/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7744 XOR2X1_7/Y XOR2X1_7/A XOR2X1_7/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7745 XOR2X1_7/a_35_54# XOR2X1_7/a_2_6# XOR2X1_7/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7746 vdd NOR2X1_2/Y XOR2X1_7/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7747 XOR2X1_7/a_13_43# NOR2X1_2/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7748 gnd XOR2X1_7/A XOR2X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7749 XOR2X1_7/a_18_6# XOR2X1_7/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7750 XOR2X1_7/Y XOR2X1_7/a_2_6# XOR2X1_7/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7751 XOR2X1_7/a_35_6# XOR2X1_7/A XOR2X1_7/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7752 gnd NOR2X1_2/Y XOR2X1_7/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7753 XOR2X1_7/a_13_43# NOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7754 vdd NOR2X1_2/A AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=440 ps=182
M7755 AOI21X1_1/a_2_54# NOR2X1_2/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7756 INVX2_6/A NOR2X1_2/Y AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7757 AOI21X1_1/a_12_6# NOR2X1_2/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7758 INVX2_6/A NOR2X1_2/B AOI21X1_1/a_12_6# Gnd nfet w=20 l=2
+  ad=110 pd=52 as=0 ps=0
M7759 gnd NOR2X1_2/Y INVX2_6/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7760 NOR2X1_2/a_9_54# NOR2X1_2/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7761 NOR2X1_2/Y NOR2X1_2/B NOR2X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7762 NOR2X1_2/Y NOR2X1_2/A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M7763 gnd NOR2X1_2/B NOR2X1_2/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7764 vdd INVX2_5/A XNOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7765 XNOR2X1_2/a_18_54# XNOR2X1_2/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7766 AND2X2_5/A XNOR2X1_2/a_2_6# XNOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7767 XNOR2X1_2/a_35_54# INVX2_5/A AND2X2_5/A vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7768 vdd XOR2X1_9/Y XNOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7769 XNOR2X1_2/a_12_41# XOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7770 gnd INVX2_5/A XNOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7771 XNOR2X1_2/a_18_6# XNOR2X1_2/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7772 AND2X2_5/A INVX2_5/A XNOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7773 XNOR2X1_2/a_35_6# XNOR2X1_2/a_2_6# AND2X2_5/A Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7774 gnd XOR2X1_9/Y XNOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7775 XNOR2X1_2/a_12_41# XOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7776 INVX2_4/Y INVX2_4/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7777 INVX2_4/Y INVX2_4/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7778 NOR2X1_1/a_9_54# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7779 XOR2X1_2/B XOR2X1_3/B NOR2X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7780 XOR2X1_2/B INVX2_4/Y gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M7781 gnd XOR2X1_3/B XOR2X1_2/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7782 vdd INVX2_4/A XOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7783 XOR2X1_3/a_18_54# XOR2X1_3/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7784 XOR2X1_3/Y INVX2_4/A XOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7785 XOR2X1_3/a_35_54# XOR2X1_3/a_2_6# XOR2X1_3/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7786 vdd XOR2X1_3/B XOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7787 XOR2X1_3/a_13_43# XOR2X1_3/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7788 gnd INVX2_4/A XOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7789 XOR2X1_3/a_18_6# XOR2X1_3/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7790 XOR2X1_3/Y XOR2X1_3/a_2_6# XOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7791 XOR2X1_3/a_35_6# INVX2_4/A XOR2X1_3/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7792 gnd XOR2X1_3/B XOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7793 XOR2X1_3/a_13_43# XOR2X1_3/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7794 vdd XOR2X1_2/A XOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7795 XOR2X1_2/a_18_54# XOR2X1_2/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7796 XOR2X1_2/Y XOR2X1_2/A XOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7797 XOR2X1_2/a_35_54# XOR2X1_2/a_2_6# XOR2X1_2/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7798 vdd XOR2X1_2/B XOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7799 XOR2X1_2/a_13_43# XOR2X1_2/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7800 gnd XOR2X1_2/A XOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7801 XOR2X1_2/a_18_6# XOR2X1_2/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7802 XOR2X1_2/Y XOR2X1_2/a_2_6# XOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7803 XOR2X1_2/a_35_6# XOR2X1_2/A XOR2X1_2/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7804 gnd XOR2X1_2/B XOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7805 XOR2X1_2/a_13_43# XOR2X1_2/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7806 OAI21X1_3/a_9_54# OAI21X1_2/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7807 XOR2X1_2/A XOR2X1_3/Y OAI21X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7808 vdd NAND3X1_0/Y XOR2X1_2/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7809 gnd OAI21X1_2/A OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7810 OAI21X1_3/a_2_6# XOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7811 XOR2X1_2/A NAND3X1_0/Y OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7812 NAND3X1_0/Y AND2X2_4/A vdd vdd pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M7813 vdd OAI21X1_2/C NAND3X1_0/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7814 NAND3X1_0/Y XOR2X1_1/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7815 NAND3X1_0/a_9_6# AND2X2_4/A gnd Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7816 NAND3X1_0/a_14_6# OAI21X1_2/C NAND3X1_0/a_9_6# Gnd nfet w=30 l=2
+  ad=90 pd=66 as=0 ps=0
M7817 NAND3X1_0/Y XOR2X1_1/B NAND3X1_0/a_14_6# Gnd nfet w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M7818 OAI21X1_2/C OAI21X1_2/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7819 vdd XOR2X1_3/Y OAI21X1_2/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7820 NAND2X1_1/a_9_6# OAI21X1_2/A gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7821 OAI21X1_2/C XOR2X1_3/Y NAND2X1_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7822 OAI21X1_2/a_9_54# OAI21X1_2/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7823 XNOR2X1_0/A XOR2X1_3/Y OAI21X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7824 vdd OAI21X1_2/C XNOR2X1_0/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7825 gnd OAI21X1_2/A OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7826 OAI21X1_2/a_2_6# XOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7827 XNOR2X1_0/A OAI21X1_2/C OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7828 AND2X2_4/a_2_6# AND2X2_4/A vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7829 vdd XOR2X1_1/B AND2X2_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7830 AND2X2_4/Y AND2X2_4/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7831 AND2X2_4/a_9_6# AND2X2_4/A AND2X2_4/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7832 gnd XOR2X1_1/B AND2X2_4/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7833 AND2X2_4/Y AND2X2_4/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7834 vdd XNOR2X1_0/A XNOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7835 XNOR2X1_0/a_18_54# XNOR2X1_0/a_12_41# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7836 XNOR2X1_0/Y XNOR2X1_0/a_2_6# XNOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7837 XNOR2X1_0/a_35_54# XNOR2X1_0/A XNOR2X1_0/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7838 vdd AND2X2_4/Y XNOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7839 XNOR2X1_0/a_12_41# AND2X2_4/Y vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7840 gnd XNOR2X1_0/A XNOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7841 XNOR2X1_0/a_18_6# XNOR2X1_0/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7842 XNOR2X1_0/Y XNOR2X1_0/A XNOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7843 XNOR2X1_0/a_35_6# XNOR2X1_0/a_2_6# XNOR2X1_0/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7844 gnd AND2X2_4/Y XNOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7845 XNOR2X1_0/a_12_41# AND2X2_4/Y gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7846 INVX2_3/Y INVX2_3/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7847 INVX2_3/Y INVX2_3/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7848 vdd XOR2X1_0/A XOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7849 XOR2X1_0/a_18_54# XOR2X1_0/a_13_43# vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7850 XOR2X1_0/Y XOR2X1_0/A XOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M7851 XOR2X1_0/a_35_54# XOR2X1_0/a_2_6# XOR2X1_0/Y vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7852 vdd XOR2X1_0/B XOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7853 XOR2X1_0/a_13_43# XOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7854 gnd XOR2X1_0/A XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7855 XOR2X1_0/a_18_6# XOR2X1_0/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7856 XOR2X1_0/Y XOR2X1_0/a_2_6# XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M7857 XOR2X1_0/a_35_6# XOR2X1_0/A XOR2X1_0/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7858 gnd XOR2X1_0/B XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7859 XOR2X1_0/a_13_43# XOR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7860 OAI21X1_0/a_9_54# OAI21X1_0/A vdd vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M7861 XOR2X1_0/A INVX2_3/Y OAI21X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M7862 vdd NAND3X1_2/Y XOR2X1_0/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7863 gnd OAI21X1_0/A OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M7864 OAI21X1_0/a_2_6# INVX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7865 XOR2X1_0/A NAND3X1_2/Y OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7866 vdd INVX2_41/Y DFFPOSX1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7867 DFFPOSX1_6/a_17_74# INVX2_2/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7868 DFFPOSX1_6/a_22_6# INVX2_41/Y DFFPOSX1_6/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7869 DFFPOSX1_6/a_31_74# DFFPOSX1_6/a_2_6# DFFPOSX1_6/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7870 vdd DFFPOSX1_6/a_34_4# DFFPOSX1_6/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7871 DFFPOSX1_6/a_34_4# DFFPOSX1_6/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7872 DFFPOSX1_6/a_61_74# DFFPOSX1_6/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7873 DFFPOSX1_6/a_66_6# DFFPOSX1_6/a_2_6# DFFPOSX1_6/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7874 DFFPOSX1_6/a_76_84# INVX2_41/Y DFFPOSX1_6/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7875 vdd con_countWriteout[4] DFFPOSX1_6/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7876 gnd INVX2_41/Y DFFPOSX1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7877 con_countWriteout[4] DFFPOSX1_6/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7878 DFFPOSX1_6/a_17_6# INVX2_2/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7879 DFFPOSX1_6/a_22_6# DFFPOSX1_6/a_2_6# DFFPOSX1_6/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7880 DFFPOSX1_6/a_31_6# INVX2_41/Y DFFPOSX1_6/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7881 gnd DFFPOSX1_6/a_34_4# DFFPOSX1_6/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7882 DFFPOSX1_6/a_34_4# DFFPOSX1_6/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7883 DFFPOSX1_6/a_61_6# DFFPOSX1_6/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7884 DFFPOSX1_6/a_66_6# INVX2_41/Y DFFPOSX1_6/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7885 DFFPOSX1_6/a_76_6# DFFPOSX1_6/a_2_6# DFFPOSX1_6/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7886 gnd con_countWriteout[4] DFFPOSX1_6/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7887 con_countWriteout[4] DFFPOSX1_6/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7888 vdd BUFX2_5/Y DFFPOSX1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7889 DFFPOSX1_5/a_17_74# AND2X2_3/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7890 DFFPOSX1_5/a_22_6# BUFX2_5/Y DFFPOSX1_5/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7891 DFFPOSX1_5/a_31_74# DFFPOSX1_5/a_2_6# DFFPOSX1_5/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7892 vdd DFFPOSX1_5/a_34_4# DFFPOSX1_5/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7893 DFFPOSX1_5/a_34_4# DFFPOSX1_5/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7894 DFFPOSX1_5/a_61_74# DFFPOSX1_5/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7895 DFFPOSX1_5/a_66_6# DFFPOSX1_5/a_2_6# DFFPOSX1_5/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7896 DFFPOSX1_5/a_76_84# BUFX2_5/Y DFFPOSX1_5/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7897 vdd AOI22X1_3/C DFFPOSX1_5/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7898 gnd BUFX2_5/Y DFFPOSX1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7899 AOI22X1_3/C DFFPOSX1_5/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7900 DFFPOSX1_5/a_17_6# AND2X2_3/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7901 DFFPOSX1_5/a_22_6# DFFPOSX1_5/a_2_6# DFFPOSX1_5/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7902 DFFPOSX1_5/a_31_6# BUFX2_5/Y DFFPOSX1_5/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7903 gnd DFFPOSX1_5/a_34_4# DFFPOSX1_5/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7904 DFFPOSX1_5/a_34_4# DFFPOSX1_5/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7905 DFFPOSX1_5/a_61_6# DFFPOSX1_5/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7906 DFFPOSX1_5/a_66_6# BUFX2_5/Y DFFPOSX1_5/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7907 DFFPOSX1_5/a_76_6# DFFPOSX1_5/a_2_6# DFFPOSX1_5/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7908 gnd AOI22X1_3/C DFFPOSX1_5/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7909 AOI22X1_3/C DFFPOSX1_5/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7910 AND2X2_3/a_2_6# HAX1_3/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7911 vdd AND2X2_6/B AND2X2_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7912 AND2X2_3/Y AND2X2_3/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7913 AND2X2_3/a_9_6# HAX1_3/YS AND2X2_3/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7914 gnd AND2X2_6/B AND2X2_3/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7915 AND2X2_3/Y AND2X2_3/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7916 INVX2_0/Y INVX2_0/A vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7917 INVX2_0/Y INVX2_0/A gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7918 vdd INVX2_41/Y DFFPOSX1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7919 DFFPOSX1_3/a_17_74# INVX2_0/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7920 DFFPOSX1_3/a_22_6# INVX2_41/Y DFFPOSX1_3/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7921 DFFPOSX1_3/a_31_74# DFFPOSX1_3/a_2_6# DFFPOSX1_3/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7922 vdd DFFPOSX1_3/a_34_4# DFFPOSX1_3/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7923 DFFPOSX1_3/a_34_4# DFFPOSX1_3/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7924 DFFPOSX1_3/a_61_74# DFFPOSX1_3/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7925 DFFPOSX1_3/a_66_6# DFFPOSX1_3/a_2_6# DFFPOSX1_3/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7926 DFFPOSX1_3/a_76_84# INVX2_41/Y DFFPOSX1_3/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7927 vdd con_countWriteout[5] DFFPOSX1_3/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7928 gnd INVX2_41/Y DFFPOSX1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7929 con_countWriteout[5] DFFPOSX1_3/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7930 DFFPOSX1_3/a_17_6# INVX2_0/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7931 DFFPOSX1_3/a_22_6# DFFPOSX1_3/a_2_6# DFFPOSX1_3/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7932 DFFPOSX1_3/a_31_6# INVX2_41/Y DFFPOSX1_3/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7933 gnd DFFPOSX1_3/a_34_4# DFFPOSX1_3/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7934 DFFPOSX1_3/a_34_4# DFFPOSX1_3/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7935 DFFPOSX1_3/a_61_6# DFFPOSX1_3/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7936 DFFPOSX1_3/a_66_6# INVX2_41/Y DFFPOSX1_3/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7937 DFFPOSX1_3/a_76_6# DFFPOSX1_3/a_2_6# DFFPOSX1_3/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7938 gnd con_countWriteout[5] DFFPOSX1_3/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7939 con_countWriteout[5] DFFPOSX1_3/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7940 AND2X2_2/a_2_6# HAX1_2/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7941 vdd AND2X2_6/B AND2X2_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7942 AND2X2_2/Y AND2X2_2/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7943 AND2X2_2/a_9_6# HAX1_2/YS AND2X2_2/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7944 gnd AND2X2_6/B AND2X2_2/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7945 AND2X2_2/Y AND2X2_2/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7946 AND2X2_1/a_2_6# HAX1_1/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7947 vdd AND2X2_6/B AND2X2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7948 AND2X2_1/Y AND2X2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7949 AND2X2_1/a_9_6# HAX1_1/YS AND2X2_1/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7950 gnd AND2X2_6/B AND2X2_1/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7951 AND2X2_1/Y AND2X2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7952 vdd BUFX2_5/Y DFFPOSX1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7953 DFFPOSX1_2/a_17_74# AND2X2_1/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7954 DFFPOSX1_2/a_22_6# BUFX2_5/Y DFFPOSX1_2/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7955 DFFPOSX1_2/a_31_74# DFFPOSX1_2/a_2_6# DFFPOSX1_2/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7956 vdd DFFPOSX1_2/a_34_4# DFFPOSX1_2/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7957 DFFPOSX1_2/a_34_4# DFFPOSX1_2/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7958 DFFPOSX1_2/a_61_74# DFFPOSX1_2/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7959 DFFPOSX1_2/a_66_6# DFFPOSX1_2/a_2_6# DFFPOSX1_2/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7960 DFFPOSX1_2/a_76_84# BUFX2_5/Y DFFPOSX1_2/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7961 vdd AOI22X1_1/C DFFPOSX1_2/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7962 gnd BUFX2_5/Y DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7963 AOI22X1_1/C DFFPOSX1_2/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7964 DFFPOSX1_2/a_17_6# AND2X2_1/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7965 DFFPOSX1_2/a_22_6# DFFPOSX1_2/a_2_6# DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7966 DFFPOSX1_2/a_31_6# BUFX2_5/Y DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7967 gnd DFFPOSX1_2/a_34_4# DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7968 DFFPOSX1_2/a_34_4# DFFPOSX1_2/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7969 DFFPOSX1_2/a_61_6# DFFPOSX1_2/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7970 DFFPOSX1_2/a_66_6# BUFX2_5/Y DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7971 DFFPOSX1_2/a_76_6# DFFPOSX1_2/a_2_6# DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7972 gnd AOI22X1_1/C DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7973 AOI22X1_1/C DFFPOSX1_2/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7974 AND2X2_0/a_2_6# HAX1_0/YS vdd vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7975 vdd AND2X2_6/B AND2X2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7976 AND2X2_0/Y AND2X2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7977 AND2X2_0/a_9_6# HAX1_0/YS AND2X2_0/a_2_6# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=100 ps=50
M7978 gnd AND2X2_6/B AND2X2_0/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7979 AND2X2_0/Y AND2X2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7980 vdd BUFX2_5/Y DFFPOSX1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M7981 DFFPOSX1_1/a_17_74# AND2X2_0/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7982 DFFPOSX1_1/a_22_6# BUFX2_5/Y DFFPOSX1_1/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M7983 DFFPOSX1_1/a_31_74# DFFPOSX1_1/a_2_6# DFFPOSX1_1/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M7984 vdd DFFPOSX1_1/a_34_4# DFFPOSX1_1/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7985 DFFPOSX1_1/a_34_4# DFFPOSX1_1/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M7986 DFFPOSX1_1/a_61_74# DFFPOSX1_1/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M7987 DFFPOSX1_1/a_66_6# DFFPOSX1_1/a_2_6# DFFPOSX1_1/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M7988 DFFPOSX1_1/a_76_84# BUFX2_5/Y DFFPOSX1_1/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7989 vdd AOI22X1_0/C DFFPOSX1_1/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7990 gnd BUFX2_5/Y DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M7991 AOI22X1_0/C DFFPOSX1_1/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M7992 DFFPOSX1_1/a_17_6# AND2X2_0/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7993 DFFPOSX1_1/a_22_6# DFFPOSX1_1/a_2_6# DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7994 DFFPOSX1_1/a_31_6# BUFX2_5/Y DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7995 gnd DFFPOSX1_1/a_34_4# DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7996 DFFPOSX1_1/a_34_4# DFFPOSX1_1/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M7997 DFFPOSX1_1/a_61_6# DFFPOSX1_1/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M7998 DFFPOSX1_1/a_66_6# BUFX2_5/Y DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M7999 DFFPOSX1_1/a_76_6# DFFPOSX1_1/a_2_6# DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8000 gnd AOI22X1_0/C DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8001 AOI22X1_0/C DFFPOSX1_1/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M8002 vdd INVX2_41/Y DFFPOSX1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M8003 DFFPOSX1_0/a_17_74# INVX2_1/Y vdd vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M8004 DFFPOSX1_0/a_22_6# INVX2_41/Y DFFPOSX1_0/a_17_74# vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M8005 DFFPOSX1_0/a_31_74# DFFPOSX1_0/a_2_6# DFFPOSX1_0/a_22_6# vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M8006 vdd DFFPOSX1_0/a_34_4# DFFPOSX1_0/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8007 DFFPOSX1_0/a_34_4# DFFPOSX1_0/a_22_6# vdd vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M8008 DFFPOSX1_0/a_61_74# DFFPOSX1_0/a_34_4# vdd vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M8009 DFFPOSX1_0/a_66_6# DFFPOSX1_0/a_2_6# DFFPOSX1_0/a_61_74# vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M8010 DFFPOSX1_0/a_76_84# INVX2_41/Y DFFPOSX1_0/a_66_6# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8011 vdd con_countWriteout[7] DFFPOSX1_0/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8012 gnd INVX2_41/Y DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M8013 con_countWriteout[7] DFFPOSX1_0/a_66_6# vdd vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M8014 DFFPOSX1_0/a_17_6# INVX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8015 DFFPOSX1_0/a_22_6# DFFPOSX1_0/a_2_6# DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8016 DFFPOSX1_0/a_31_6# INVX2_41/Y DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8017 gnd DFFPOSX1_0/a_34_4# DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8018 DFFPOSX1_0/a_34_4# DFFPOSX1_0/a_22_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M8019 DFFPOSX1_0/a_61_6# DFFPOSX1_0/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8020 DFFPOSX1_0/a_66_6# INVX2_41/Y DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M8021 DFFPOSX1_0/a_76_6# DFFPOSX1_0/a_2_6# DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M8022 gnd con_countWriteout[7] DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8023 con_countWriteout[7] DFFPOSX1_0/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 vdd XNOR2X1_23/a_2_6# 2.29fF
C1 vdd OAI21X1_87/C 6.26fF
C2 vdd con_restart 59.61fF
C3 vdd INVX2_59/Y 10.04fF
C4 vdd DFFPOSX1_7/a_2_6# 5.17fF
C5 out_MuxData[12] out_MuxData[13] 2.57fF
C6 vdd OAI21X1_59/B 3.53fF
C7 vdd DFFPOSX1_91/a_2_6# 5.17fF
C8 out_MuxData[13] gnd 18.59fF
C9 AOI22X1_26/a_2_54# vdd 2.85fF
C10 DFFPOSX1_64/a_22_6# vdd 2.55fF
C11 XNOR2X1_34/a_2_6# OAI21X1_58/Y 2.10fF
C12 vdd DFFPOSX1_74/a_34_4# 2.60fF
C13 vdd XOR2X1_4/Y 4.16fF
C14 vdd XOR2X1_47/Y 5.86fF
C15 vdd XOR2X1_17/B 41.04fF
C16 vdd XOR2X1_43/Y 3.30fF
C17 out_MuxData[10] INVX2_17/Y 2.95fF
C18 con_readData gnd 12.32fF
C19 vdd XOR2X1_89/a_13_43# 2.11fF
C20 out_MemBData[4] gnd 4.17fF
C21 INVX2_109/Y vdd 8.58fF
C22 vdd DFFPOSX1_76/a_34_4# 2.60fF
C23 vdd AOI22X1_23/a_2_54# 2.85fF
C24 vdd XOR2X1_81/a_2_6# 2.07fF
C25 gnd INVX2_17/Y 15.32fF
C26 vdd DFFPOSX1_24/a_2_6# 5.17fF
C27 vdd AOI22X1_1/C 2.68fF
C28 OAI21X1_68/B vdd 8.31fF
C29 INVX2_126/A con_count[0] 2.42fF
C30 XOR2X1_90/A gnd 2.13fF
C31 out_MuxData[1] out_MuxData[0] 4.19fF
C32 vdd INVX2_26/A 25.09fF
C33 XNOR2X1_58/A AND2X2_38/Y 3.16fF
C34 XOR2X1_59/a_13_43# vdd 2.11fF
C35 vdd HAX1_10/YS 6.25fF
C36 vdd XOR2X1_90/a_13_43# 2.11fF
C37 AND2X2_17/Y gnd 2.60fF
C38 vdd DFFPOSX1_90/a_34_4# 2.60fF
C39 out_MuxData[7] INVX2_28/Y 2.12fF
C40 vdd DFFPOSX1_0/a_22_6# 2.55fF
C41 INVX2_50/Y gnd 3.23fF
C42 vdd XOR2X1_55/A 7.07fF
C43 AOI22X1_41/Y AOI22X1_41/a_2_54# 2.15fF
C44 AND2X2_39/B NOR2X1_46/B 2.31fF
C45 vdd DFFPOSX1_39/a_22_6# 2.55fF
C46 in_clkb DFFPOSX1_31/a_22_6# 2.18fF
C47 vdd OAI21X1_47/C 4.62fF
C48 vdd OAI21X1_56/A 8.91fF
C49 vdd OAI21X1_83/Y 4.39fF
C50 vdd DFFPOSX1_32/a_34_4# 2.60fF
C51 vdd HAX1_2/YS 3.00fF
C52 vdd AND2X2_1/Y 3.15fF
C53 vdd NAND3X1_15/Y 6.91fF
C54 vdd AOI22X1_97/a_2_54# 2.85fF
C55 vdd XOR2X1_87/Y 2.82fF
C56 AND2X2_36/A DFFPOSX1_71/a_34_4# 2.39fF
C57 out_MuxData[1] XOR2X1_52/a_2_6# 2.42fF
C58 vdd DFFPOSX1_29/a_34_4# 2.60fF
C59 vdd OAI21X1_60/C 6.91fF
C60 vdd NAND3X1_8/B 3.89fF
C61 BUFX2_9/Y gnd 22.91fF
C62 vdd XOR2X1_40/a_2_6# 2.07fF
C63 DFFPOSX1_2/a_22_6# vdd 2.55fF
C64 XOR2X1_17/a_2_6# vdd 2.07fF
C65 XOR2X1_65/a_13_43# out_MuxData[10] 2.33fF
C66 INVX2_41/Y DFFPOSX1_45/a_22_6# 2.18fF
C67 vdd XOR2X1_31/a_13_43# 2.04fF
C68 vdd XOR2X1_55/a_13_43# 2.11fF
C69 AOI22X1_18/a_2_54# vdd 2.85fF
C70 XOR2X1_87/B vdd 12.96fF
C71 in_inp vdd 8.53fF
C72 vdd DFFPOSX1_32/a_2_6# 5.17fF
C73 vdd AOI22X1_32/a_2_54# 2.85fF
C74 vdd AOI22X1_58/a_2_54# 2.85fF
C75 out_MemBData[10] gnd 2.89fF
C76 vdd AOI22X1_30/Y 8.58fF
C77 vdd XNOR2X1_36/a_2_6# 2.29fF
C78 INVX2_86/A out_MuxData[13] 2.64fF
C79 vdd DFFPOSX1_42/a_2_6# 5.17fF
C80 vdd INVX2_87/Y 36.61fF
C81 BUFX2_9/Y DFFPOSX1_16/a_22_6# 2.16fF
C82 XOR2X1_13/a_2_6# vdd 2.07fF
C83 AND2X2_27/Y vdd 3.11fF
C84 DFFPOSX1_35/a_22_6# vdd 2.55fF
C85 vdd XOR2X1_75/a_13_43# 2.11fF
C86 vdd AOI22X1_79/C 2.68fF
C87 vdd DFFPOSX1_78/a_34_4# 2.60fF
C88 DFFPOSX1_38/a_2_6# vdd 5.17fF
C89 XOR2X1_13/Y vdd 4.55fF
C90 AOI22X1_69/a_2_54# vdd 2.85fF
C91 vdd out_MemBData[11] 12.46fF
C92 vdd out_MuxData[8] 56.29fF
C93 vdd out_MemBData[9] 15.37fF
C94 vdd OAI21X1_62/Y 2.88fF
C95 AOI22X1_19/C AND2X2_6/B 2.47fF
C96 vdd DFFPOSX1_1/a_34_4# 2.60fF
C97 INVX2_104/Y vdd 33.49fF
C98 XOR2X1_35/Y vdd 4.88fF
C99 XOR2X1_71/a_2_6# vdd 2.07fF
C100 vdd INVX2_84/Y 25.71fF
C101 vdd INVX2_120/A 7.11fF
C102 NOR2X1_12/A vdd 6.02fF
C103 INVX2_41/Y DFFPOSX1_7/a_2_6# 3.07fF
C104 vdd AOI22X1_62/B 8.64fF
C105 vdd DFFPOSX1_22/a_22_6# 2.55fF
C106 vdd AOI22X1_33/a_2_54# 2.85fF
C107 vdd INVX2_9/A 2.94fF
C108 vdd XOR2X1_64/B 2.10fF
C109 vdd NOR2X1_0/B 4.85fF
C110 out_MuxData[12] XOR2X1_9/a_2_6# 2.34fF
C111 vdd AND2X2_39/Y 30.68fF
C112 vdd con_countWriteout[3] 11.66fF
C113 vdd DFFPOSX1_28/a_34_4# 2.60fF
C114 XOR2X1_36/B out_MuxData[5] 2.10fF
C115 INVX2_126/A INVX2_72/Y 2.42fF
C116 AND2X2_5/A gnd 6.34fF
C117 vdd XOR2X1_79/a_13_43# 2.11fF
C118 vdd OAI21X1_78/B 3.40fF
C119 vdd con_count[4] 11.81fF
C120 vdd DFFPOSX1_98/a_22_6# 2.55fF
C121 XOR2X1_70/a_2_6# out_MuxData[0] 2.42fF
C122 XOR2X1_26/a_13_43# AND2X2_14/A 2.06fF
C123 XOR2X1_55/B out_MuxData[2] 2.13fF
C124 vdd AOI22X1_36/a_2_54# 2.85fF
C125 vdd INVX2_131/Y 4.45fF
C126 vdd XNOR2X1_57/Y 2.95fF
C127 XNOR2X1_40/a_2_6# vdd 2.29fF
C128 out_MuxData[1] OAI22X1_6/C 2.72fF
C129 DFFPOSX1_71/a_22_6# vdd 2.55fF
C130 vdd XOR2X1_49/A 5.09fF
C131 vdd INVX2_128/A 5.67fF
C132 vdd INVX2_48/A 2.44fF
C133 vdd XOR2X1_48/a_13_43# 2.11fF
C134 vdd XOR2X1_57/a_2_6# 2.07fF
C135 vdd BUFX2_8/a_2_6# 2.41fF
C136 AND2X2_41/A XOR2X1_91/a_13_43# 2.18fF
C137 vdd XNOR2X1_18/a_2_6# 2.29fF
C138 XNOR2X1_42/a_2_6# vdd 2.29fF
C139 XOR2X1_69/a_2_6# vdd 2.07fF
C140 INVX2_16/Y INVX2_17/Y 2.12fF
C141 vdd NAND2X1_17/B 3.70fF
C142 vdd DFFPOSX1_81/a_34_4# 2.60fF
C143 DFFPOSX1_66/a_34_4# vdd 2.60fF
C144 INVX2_130/A gnd 2.50fF
C145 vdd AOI22X1_81/a_2_54# 2.85fF
C146 vdd NAND3X1_2/B 8.47fF
C147 vdd NAND2X1_42/Y 4.61fF
C148 vdd AOI22X1_83/a_2_54# 2.85fF
C149 vdd INVX2_22/Y 8.17fF
C150 INVX2_83/Y out_MuxData[4] 2.08fF
C151 vdd DFFPOSX1_93/a_2_6# 5.17fF
C152 INVX2_60/Y OR2X2_0/Y 3.03fF
C153 INVX2_11/A INVX2_36/A 2.00fF
C154 AND2X2_24/Y XNOR2X1_34/a_12_41# 2.64fF
C155 AND2X2_21/A vdd 4.29fF
C156 DFFPOSX1_61/a_34_4# vdd 2.60fF
C157 XOR2X1_24/Y vdd 11.93fF
C158 vdd AND2X2_15/Y 4.64fF
C159 DFFPOSX1_67/a_2_6# vdd 5.17fF
C160 vdd AOI22X1_48/Y 4.12fF
C161 vdd XOR2X1_4/a_13_43# 2.11fF
C162 vdd XNOR2X1_48/a_2_6# 2.29fF
C163 vdd NOR2X1_35/Y 12.54fF
C164 vdd INVX2_20/Y 4.27fF
C165 out_MuxData[1] XOR2X1_51/Y 2.01fF
C166 OR2X1_2/Y vdd 6.07fF
C167 XOR2X1_68/B vdd 6.26fF
C168 con_loadData vdd 4.64fF
C169 vdd HAX1_0/a_2_74# 3.67fF
C170 vdd INVX2_134/Y 20.47fF
C171 vdd NAND3X1_16/B 14.44fF
C172 vdd DFFPOSX1_21/a_2_6# 5.17fF
C173 XOR2X1_51/a_2_6# vdd 2.07fF
C174 vdd XNOR2X1_7/Y 3.30fF
C175 vdd DFFPOSX1_33/a_22_6# 2.55fF
C176 NAND2X1_4/Y NAND2X1_4/B 4.36fF
C177 vdd BUFX2_0/A 3.53fF
C178 vdd OAI21X1_76/C 4.62fF
C179 out_MuxData[7] out_MuxData[13] 3.92fF
C180 vdd DFFPOSX1_51/a_22_6# 2.55fF
C181 NOR2X1_17/A NOR2X1_17/B 2.11fF
C182 INVX2_11/A INVX2_1/A 2.61fF
C183 con_countWriteout[6] vdd 7.02fF
C184 DFFPOSX1_64/a_34_4# vdd 2.60fF
C185 vdd HAX1_8/YS 3.58fF
C186 vdd AOI22X1_61/a_2_54# 2.85fF
C187 XOR2X1_41/a_2_6# vdd 2.07fF
C188 AOI22X1_67/C vdd 2.68fF
C189 vdd DFFPOSX1_86/a_22_6# 2.55fF
C190 vdd BUFX2_0/a_2_6# 2.41fF
C191 INVX2_16/Y NOR2X1_8/Y 2.01fF
C192 AOI22X1_76/a_2_54# vdd 2.85fF
C193 XOR2X1_50/A vdd 4.97fF
C194 INVX2_91/Y vdd 5.81fF
C195 vdd OAI21X1_60/Y 4.65fF
C196 AND2X2_29/a_2_6# INVX2_72/Y 2.76fF
C197 vdd NAND3X1_4/Y 5.91fF
C198 XOR2X1_88/B XOR2X1_88/a_13_43# 2.64fF
C199 vdd NAND2X1_4/B 5.75fF
C200 vdd XOR2X1_54/a_2_6# 2.07fF
C201 vdd HAX1_1/B 4.91fF
C202 vdd XOR2X1_58/a_2_6# 2.07fF
C203 vdd INVX2_57/Y 7.05fF
C204 vdd NAND3X1_25/Y 5.83fF
C205 vdd AOI22X1_38/A 6.21fF
C206 BUFX2_10/Y DFFPOSX1_61/a_22_6# 2.18fF
C207 AOI22X1_48/D INVX2_94/Y 2.02fF
C208 XOR2X1_1/B vdd 6.33fF
C209 DFFPOSX1_58/a_22_6# vdd 2.55fF
C210 out_MuxData[7] INVX2_17/Y 2.70fF
C211 vdd DFFPOSX1_76/a_2_6# 5.17fF
C212 XOR2X1_66/a_13_43# out_MuxData[10] 2.64fF
C213 INVX2_126/A gnd 2.79fF
C214 vdd XOR2X1_61/a_13_43# 2.11fF
C215 INVX2_39/A out_MuxData[4] 3.26fF
C216 INVX2_5/A gnd 14.84fF
C217 vdd DFFPOSX1_21/a_22_6# 2.55fF
C218 INVX2_52/A gnd 2.04fF
C219 out_MuxData[2] out_MuxData[10] 3.30fF
C220 NAND3X1_6/Y gnd 2.50fF
C221 XOR2X1_74/a_2_6# vdd 2.07fF
C222 INVX2_92/Y BUFX2_5/Y 2.06fF
C223 XOR2X1_9/B vdd 2.83fF
C224 vdd HAX1_0/YS 3.00fF
C225 vdd XNOR2X1_13/a_2_6# 2.29fF
C226 out_MuxData[12] out_MuxData[2] 2.54fF
C227 vdd INVX2_99/Y 24.25fF
C228 vdd XOR2X1_44/a_2_6# 2.07fF
C229 out_MuxData[2] gnd 21.78fF
C230 vdd HAX1_4/YS 3.00fF
C231 vdd XOR2X1_5/A 2.72fF
C232 vdd XOR2X1_49/a_2_6# 2.07fF
C233 NOR2X1_29/A XNOR2X1_41/a_12_41# 3.84fF
C234 out_state[2] gnd 4.00fF
C235 NOR2X1_31/Y vdd 18.27fF
C236 vdd DFFPOSX1_72/a_22_6# 2.55fF
C237 vdd AOI22X1_5/a_2_54# 2.85fF
C238 INVX2_28/Y XOR2X1_39/a_13_43# 2.64fF
C239 vdd INVX2_8/Y 6.42fF
C240 vdd XOR2X1_3/Y 4.52fF
C241 vdd DFFPOSX1_83/a_22_6# 2.55fF
C242 vdd NOR2X1_17/B 2.94fF
C243 vdd XNOR2X1_1/a_2_6# 2.29fF
C244 gnd OR2X2_0/Y 7.36fF
C245 AOI21X1_7/B vdd 11.57fF
C246 AND2X2_19/Y OR2X2_0/Y 2.88fF
C247 XNOR2X1_31/a_2_6# vdd 2.29fF
C248 out_MemBData[3] gnd 2.36fF
C249 vdd DFFPOSX1_20/a_2_6# 5.17fF
C250 vdd AOI22X1_53/a_2_54# 2.85fF
C251 vdd NAND3X1_12/Y 5.60fF
C252 vdd INVX2_105/Y 6.36fF
C253 XOR2X1_69/A XOR2X1_69/B 2.58fF
C254 vdd AND2X2_9/B 9.22fF
C255 vdd AOI22X1_25/a_2_54# 2.85fF
C256 vdd DFFPOSX1_31/a_2_6# 5.17fF
C257 vdd DFFPOSX1_52/a_2_6# 5.17fF
C258 vdd XOR2X1_53/a_13_43# 2.11fF
C259 DFFPOSX1_36/a_22_6# vdd 2.55fF
C260 out_MuxData[1] gnd 10.77fF
C261 vdd out_temp_addNum[1] 3.83fF
C262 XNOR2X1_19/a_2_6# XNOR2X1_19/A 2.79fF
C263 NAND3X1_8/B INVX2_27/Y 2.12fF
C264 vdd HAX1_11/a_2_74# 3.67fF
C265 vdd INVX2_124/A 2.64fF
C266 out_MuxData[12] out_MuxData[5] 2.75fF
C267 vdd DFFPOSX1_44/a_22_6# 2.55fF
C268 vdd XNOR2X1_34/a_2_6# 2.29fF
C269 gnd out_MuxData[5] 12.33fF
C270 AOI22X1_49/a_2_54# vdd 2.85fF
C271 out_MuxData[4] out_MuxData[5] 4.74fF
C272 AOI22X1_62/a_2_54# vdd 2.85fF
C273 vdd DFFPOSX1_73/a_22_6# 2.55fF
C274 AND2X2_23/Y vdd 5.37fF
C275 vdd AOI22X1_29/C 2.68fF
C276 NAND3X1_27/Y vdd 7.93fF
C277 XOR2X1_13/Y AND2X2_8/a_2_6# 2.15fF
C278 vdd XNOR2X1_19/A 3.60fF
C279 vdd OAI21X1_59/C 8.63fF
C280 vdd XOR2X1_40/a_13_43# 2.11fF
C281 vdd XOR2X1_34/Y 2.94fF
C282 gnd BUFX2_11/Y 35.84fF
C283 INVX2_25/Y gnd 20.12fF
C284 out_MuxData[9] XOR2X1_69/B 3.63fF
C285 vdd DFFPOSX1_53/a_2_6# 5.17fF
C286 XOR2X1_71/a_13_43# vdd 2.11fF
C287 vdd DFFPOSX1_60/a_34_4# 2.60fF
C288 vdd AOI22X1_84/a_2_54# 2.85fF
C289 vdd NOR2X1_28/B 2.82fF
C290 vdd out_MemBData[14] 27.91fF
C291 vdd XOR2X1_91/A 6.26fF
C292 out_state[2] out_state[1] 2.05fF
C293 INVX2_43/Y gnd 23.57fF
C294 DFFPOSX1_84/a_22_6# BUFX2_11/Y 2.18fF
C295 vdd AND2X2_3/Y 2.74fF
C296 XOR2X1_6/A XNOR2X1_9/A 2.09fF
C297 out_MuxData[1] XOR2X1_81/A 2.22fF
C298 DFFPOSX1_56/a_2_6# vdd 5.17fF
C299 INVX2_62/Y gnd 11.30fF
C300 out_MuxData[9] XNOR2X1_33/a_2_6# 2.35fF
C301 DFFPOSX1_41/a_34_4# vdd 2.60fF
C302 XOR2X1_62/Y vdd 3.97fF
C303 vdd XNOR2X1_53/a_2_6# 2.29fF
C304 vdd con_count[5] 10.01fF
C305 vdd INVX2_42/Y 3.36fF
C306 vdd AND2X2_14/Y 5.40fF
C307 vdd AOI22X1_14/a_2_54# 2.85fF
C308 vdd OAI21X1_38/Y 3.55fF
C309 vdd AOI22X1_54/a_2_54# 2.85fF
C310 vdd DFFPOSX1_46/a_2_6# 5.17fF
C311 vdd AND2X2_4/A 4.96fF
C312 XOR2X1_67/a_2_6# vdd 2.07fF
C313 XOR2X1_72/a_13_43# vdd 2.11fF
C314 out_MuxData[7] XOR2X1_42/a_13_43# 2.29fF
C315 DFFPOSX1_71/a_34_4# vdd 2.60fF
C316 XOR2X1_53/Y XNOR2X1_35/a_12_41# 3.65fF
C317 vdd INVX2_54/Y 2.19fF
C318 vdd NOR2X1_39/A 5.12fF
C319 DFFPOSX1_70/a_22_6# vdd 2.55fF
C320 vdd INVX2_28/Y 35.01fF
C321 out_MuxData[7] XOR2X1_28/a_2_6# 2.60fF
C322 XOR2X1_54/A vdd 5.39fF
C323 vdd XNOR2X1_3/Y 5.00fF
C324 vdd INVX2_63/A 2.44fF
C325 XNOR2X1_7/A XNOR2X1_7/Y 2.04fF
C326 vdd XOR2X1_37/a_2_6# 2.07fF
C327 vdd OAI21X1_30/C 6.76fF
C328 DFFPOSX1_43/a_34_4# BUFX2_5/Y 2.36fF
C329 vdd AND2X2_18/B 8.79fF
C330 INVX2_15/Y vdd 5.05fF
C331 XOR2X1_29/Y vdd 8.22fF
C332 XOR2X1_69/a_13_43# vdd 2.11fF
C333 vdd XOR2X1_77/Y 4.52fF
C334 XNOR2X1_43/a_2_6# vdd 2.29fF
C335 vdd DFFPOSX1_88/a_34_4# 2.60fF
C336 DFFPOSX1_66/a_2_6# vdd 5.17fF
C337 vdd DFFPOSX1_45/a_34_4# 2.60fF
C338 vdd XOR2X1_50/a_2_6# 2.07fF
C339 XOR2X1_30/a_2_6# OAI22X1_6/C 2.32fF
C340 vdd DFFPOSX1_20/a_34_4# 2.60fF
C341 out_MemBData[5] gnd 5.53fF
C342 vdd AOI21X1_2/Y 9.76fF
C343 XNOR2X1_14/a_12_41# INVX2_39/A 2.64fF
C344 vdd BUFX2_5/a_2_6# 2.41fF
C345 vdd AND2X2_35/Y 4.60fF
C346 vdd AOI22X1_22/a_2_54# 2.85fF
C347 INVX2_86/A out_MuxData[1] 2.36fF
C348 AOI22X1_41/Y vdd 16.68fF
C349 DFFPOSX1_55/a_22_6# vdd 2.55fF
C350 vdd HAX1_8/a_2_74# 3.67fF
C351 vdd OAI21X1_71/C 3.16fF
C352 AOI22X1_28/a_2_54# vdd 2.85fF
C353 OAI21X1_65/Y vdd 3.22fF
C354 vdd DFFPOSX1_48/a_2_6# 5.17fF
C355 vdd DFFPOSX1_18/a_2_6# 5.17fF
C356 vdd AND2X2_18/A 10.17fF
C357 vdd DFFPOSX1_15/a_22_6# 2.55fF
C358 XOR2X1_87/B INVX2_86/Y 2.09fF
C359 vdd NAND2X1_11/Y 5.64fF
C360 vdd XOR2X1_14/B 2.92fF
C361 vdd AND2X2_6/B 28.55fF
C362 XOR2X1_43/a_2_6# vdd 2.07fF
C363 INVX2_55/A vdd 5.08fF
C364 vdd NAND3X1_22/Y 5.91fF
C365 XOR2X1_41/a_13_43# vdd 2.11fF
C366 vdd NAND2X1_7/A 4.82fF
C367 con_count[1] BUFX2_9/Y 4.15fF
C368 XOR2X1_62/B out_MuxData[10] 2.48fF
C369 vdd OAI21X1_52/C 19.12fF
C370 vdd XOR2X1_85/B 6.47fF
C371 vdd HAX1_4/B 8.52fF
C372 INVX2_43/Y DFFPOSX1_24/a_22_6# 2.03fF
C373 XOR2X1_80/a_13_43# XOR2X1_69/B 2.87fF
C374 XOR2X1_6/A vdd 3.32fF
C375 BUFX2_10/Y BUFX2_11/Y 5.44fF
C376 vdd HAX1_13/a_2_74# 3.67fF
C377 AND2X2_9/A AND2X2_9/B 2.84fF
C378 vdd XOR2X1_42/a_2_6# 2.07fF
C379 vdd AND2X2_40/A 7.75fF
C380 XOR2X1_88/a_2_6# XOR2X1_88/A 2.57fF
C381 XNOR2X1_41/Y XOR2X1_69/B 2.52fF
C382 INVX2_4/A NAND2X1_5/Y 2.33fF
C383 OAI21X1_0/A AOI22X1_12/a_2_54# 2.12fF
C384 DFFPOSX1_52/a_34_4# out_MuxData[4] 2.29fF
C385 INVX2_41/Y AOI22X1_29/C 3.26fF
C386 vdd XNOR2X1_37/a_2_6# 2.29fF
C387 OAI21X1_2/C vdd 4.41fF
C388 vdd XOR2X1_83/a_13_43# 2.11fF
C389 XOR2X1_70/B vdd 5.33fF
C390 out_MuxData[7] INVX2_5/A 2.00fF
C391 vdd DFFPOSX1_16/a_34_4# 2.60fF
C392 vdd DFFPOSX1_10/a_22_6# 2.55fF
C393 vdd OAI21X1_85/C 5.04fF
C394 vdd XOR2X1_81/a_13_43# 2.11fF
C395 vdd HAX1_13/YS 5.88fF
C396 vdd XOR2X1_3/a_13_43# 2.11fF
C397 vdd DFFPOSX1_9/a_34_4# 2.60fF
C398 NOR2X1_45/A out_MuxData[4] 2.36fF
C399 out_MuxData[10] out_MuxData[0] 2.05fF
C400 AND2X2_13/Y out_MuxData[5] 2.03fF
C401 con_countWriteout[0] gnd 3.15fF
C402 XOR2X1_74/a_13_43# vdd 2.11fF
C403 XNOR2X1_32/a_2_6# vdd 2.29fF
C404 con_count[6] gnd 5.58fF
C405 vdd INVX2_52/Y 6.80fF
C406 XOR2X1_19/Y vdd 3.30fF
C407 HAX1_7/YC vdd 6.84fF
C408 vdd INVX2_126/Y 18.05fF
C409 vdd XOR2X1_32/Y 5.50fF
C410 NOR2X1_49/B gnd 9.29fF
C411 gnd out_MuxData[0] 19.95fF
C412 vdd DFFPOSX1_90/a_2_6# 5.17fF
C413 vdd INVX2_21/Y 9.41fF
C414 vdd con_countWriteout[7] 7.90fF
C415 out_MuxData[4] out_MuxData[0] 2.56fF
C416 DFFPOSX1_12/a_34_4# vdd 2.60fF
C417 HAX1_7/a_2_74# vdd 3.67fF
C418 INVX2_93/Y AND2X2_13/A 2.01fF
C419 XOR2X1_66/a_2_6# vdd 2.07fF
C420 vdd DFFPOSX1_72/a_34_4# 2.60fF
C421 vdd XOR2X1_54/B 3.22fF
C422 con_count[2] gnd 2.65fF
C423 vdd INVX2_24/Y 6.14fF
C424 out_MuxData[1] out_MuxData[6] 2.16fF
C425 vdd AOI22X1_43/a_2_54# 2.85fF
C426 vdd AND2X2_32/Y 4.26fF
C427 DFFPOSX1_51/a_2_6# BUFX2_5/Y 2.23fF
C428 vdd DFFPOSX1_29/a_2_6# 5.17fF
C429 vdd XOR2X1_8/a_13_43# 2.11fF
C430 vdd AOI22X1_19/a_2_54# 2.85fF
C431 vdd INVX2_69/Y 5.39fF
C432 gnd NOR2X1_41/B 5.53fF
C433 INVX2_104/Y con_restart 3.23fF
C434 AOI22X1_73/a_2_54# vdd 2.85fF
C435 vdd XOR2X1_9/a_13_43# 2.11fF
C436 INVX2_32/Y vdd 5.39fF
C437 out_MuxData[8] XOR2X1_17/B 2.85fF
C438 vdd DFFPOSX1_87/a_2_6# 5.17fF
C439 DFFPOSX1_60/a_22_6# vdd 2.55fF
C440 vdd AOI22X1_47/a_2_54# 2.85fF
C441 vdd XOR2X1_46/a_13_43# 2.11fF
C442 vdd DFFPOSX1_92/a_22_6# 2.55fF
C443 vdd in_clka 14.61fF
C444 vdd XOR2X1_69/B 42.53fF
C445 vdd AOI22X1_66/a_2_54# 2.85fF
C446 NOR2X1_12/A XOR2X1_43/Y 2.10fF
C447 vdd OAI21X1_71/Y 3.92fF
C448 AOI22X1_77/a_2_54# vdd 2.85fF
C449 XOR2X1_70/Y vdd 2.50fF
C450 vdd XNOR2X1_27/Y 7.31fF
C451 vdd INVX2_0/Y 2.39fF
C452 vdd XNOR2X1_47/a_2_6# 2.29fF
C453 vdd AOI22X1_50/B 4.32fF
C454 vdd HAX1_11/B 3.34fF
C455 vdd AOI22X1_87/a_2_54# 2.85fF
C456 vdd INVX2_79/Y 6.00fF
C457 vdd OAI21X1_78/C 7.27fF
C458 vdd AOI22X1_12/a_2_54# 2.85fF
C459 vdd DFFPOSX1_43/a_22_6# 2.55fF
C460 NOR2X1_27/A out_MuxData[13] 2.00fF
C461 vdd NOR2X1_8/B 7.15fF
C462 vdd out_MuxData[13] 62.37fF
C463 XOR2X1_12/a_13_43# vdd 2.11fF
C464 DFFPOSX1_35/a_34_4# vdd 2.60fF
C465 DFFPOSX1_65/a_22_6# vdd 2.55fF
C466 INVX2_56/Y vdd 18.99fF
C467 out_MemBData[1] gnd 5.23fF
C468 DFFPOSX1_14/a_2_6# vdd 5.17fF
C469 vdd XOR2X1_46/Y 3.65fF
C470 con_count[0] gnd 10.49fF
C471 vdd con_writeData 19.11fF
C472 vdd HAX1_1/a_2_74# 3.67fF
C473 vdd XNOR2X1_33/a_2_6# 2.29fF
C474 vdd con_readData 12.34fF
C475 vdd XNOR2X1_58/A 4.72fF
C476 vdd DFFPOSX1_52/a_22_6# 2.55fF
C477 INVX2_41/Y AND2X2_6/B 2.62fF
C478 vdd DFFPOSX1_96/a_34_4# 2.60fF
C479 out_MuxData[3] out_MuxData[2] 2.05fF
C480 DFFPOSX1_20/a_22_6# vdd 2.55fF
C481 DFFPOSX1_5/a_34_4# vdd 2.60fF
C482 out_MemBData[4] vdd 18.50fF
C483 DFFPOSX1_7/a_34_4# vdd 2.60fF
C484 out_MemBData[13] gnd 3.36fF
C485 AOI22X1_72/a_2_54# vdd 2.85fF
C486 OAI22X1_10/Y INVX2_99/Y 2.65fF
C487 vdd INVX2_70/Y 10.42fF
C488 vdd INVX2_17/Y 41.54fF
C489 XOR2X1_35/a_2_6# out_MuxData[5] 3.60fF
C490 vdd XOR2X1_19/a_13_43# 2.11fF
C491 vdd DFFPOSX1_28/a_2_6# 5.17fF
C492 vdd AOI22X1_30/a_2_54# 2.85fF
C493 OAI21X1_50/A out_MuxData[13] 2.74fF
C494 out_MuxData[4] XOR2X1_36/a_2_6# 2.03fF
C495 INVX2_26/Y vdd 36.05fF
C496 XOR2X1_90/A vdd 11.73fF
C497 in_clkb gnd 16.98fF
C498 vdd AND2X2_17/Y 24.58fF
C499 vdd OAI22X1_19/Y 3.62fF
C500 XOR2X1_0/a_13_43# XOR2X1_0/Y 2.02fF
C501 XNOR2X1_44/a_2_6# XOR2X1_69/A 2.10fF
C502 INVX2_41/Y DFFPOSX1_10/a_22_6# 2.47fF
C503 DFFPOSX1_71/a_2_6# vdd 5.17fF
C504 out_MuxData[9] NAND2X1_28/Y 3.04fF
C505 vdd INVX2_50/Y 17.21fF
C506 XOR2X1_75/a_13_43# INVX2_87/Y 3.82fF
C507 OAI22X1_6/C OAI21X1_40/A 2.22fF
C508 vdd NOR2X1_28/Y 5.83fF
C509 INVX2_96/A vdd 3.14fF
C510 out_MuxData[8] INVX2_87/Y 2.73fF
C511 OAI22X1_6/C gnd 12.09fF
C512 vdd NAND2X1_9/A 2.73fF
C513 vdd in_wai 14.21fF
C514 vdd OAI21X1_6/B 8.46fF
C515 vdd XOR2X1_91/a_2_6# 2.07fF
C516 XOR2X1_3/Y NAND3X1_0/Y 2.04fF
C517 vdd XOR2X1_39/a_2_6# 2.07fF
C518 BUFX2_10/Y DFFPOSX1_70/a_2_6# 2.02fF
C519 AOI22X1_55/D vdd 4.36fF
C520 INVX2_67/Y INVX2_92/Y 3.73fF
C521 NAND3X1_1/Y vdd 4.86fF
C522 DFFPOSX1_56/a_22_6# vdd 2.55fF
C523 INVX2_53/Y INVX2_43/Y 2.69fF
C524 vdd DFFPOSX1_81/a_2_6# 5.17fF
C525 INVX2_93/Y INVX2_49/A 2.22fF
C526 vdd DFFPOSX1_88/a_2_6# 5.17fF
C527 OAI21X1_67/C vdd 7.13fF
C528 vdd BUFX2_9/Y 70.39fF
C529 vdd AND2X2_39/B 3.85fF
C530 vdd XOR2X1_22/A 2.53fF
C531 NOR2X1_15/B AND2X2_20/Y 2.46fF
C532 vdd XOR2X1_78/a_13_43# 2.11fF
C533 vdd XOR2X1_83/B 2.33fF
C534 vdd DFFPOSX1_12/a_2_6# 5.17fF
C535 AND2X2_28/B vdd 13.99fF
C536 DFFPOSX1_61/a_2_6# vdd 5.17fF
C537 DFFPOSX1_23/a_22_6# vdd 2.55fF
C538 vdd XOR2X1_7/a_2_6# 2.07fF
C539 vdd DFFPOSX1_86/a_2_6# 5.17fF
C540 vdd XOR2X1_33/A 2.67fF
C541 DFFPOSX1_7/a_22_6# vdd 2.55fF
C542 vdd DFFPOSX1_1/a_22_6# 2.55fF
C543 vdd out_MemBData[10] 16.20fF
C544 vdd NOR2X1_23/Y 3.37fF
C545 vdd XOR2X1_43/B 7.02fF
C546 AND2X2_3/Y con_countWriteout[2] 3.16fF
C547 INVX2_107/A vdd 2.59fF
C548 vdd XOR2X1_65/a_13_43# 2.11fF
C549 vdd HAX1_12/a_2_74# 3.67fF
C550 vdd XOR2X1_65/Y 6.33fF
C551 INVX2_72/Y gnd 2.31fF
C552 vdd DFFPOSX1_1/a_2_6# 5.17fF
C553 con_countWriteout[5] gnd 5.14fF
C554 vdd NAND3X1_7/Y 10.17fF
C555 vdd DFFPOSX1_49/a_22_6# 2.55fF
C556 vdd HAX1_0/YC 3.85fF
C557 vdd AOI22X1_4/a_2_54# 2.85fF
C558 vdd INVX2_7/Y 2.46fF
C559 vdd OAI21X1_61/Y 4.51fF
C560 vdd XOR2X1_50/B 4.76fF
C561 vdd XNOR2X1_58/a_2_6# 2.29fF
C562 vdd out_MemBData[15] 11.85fF
C563 vdd XOR2X1_54/Y 2.89fF
C564 NAND3X1_8/C vdd 7.18fF
C565 DFFPOSX1_64/a_2_6# vdd 5.17fF
C566 DFFPOSX1_61/a_22_6# vdd 2.55fF
C567 out_MemBData[12] gnd 2.26fF
C568 vdd XOR2X1_47/a_13_43# 2.11fF
C569 XOR2X1_71/Y vdd 4.79fF
C570 INVX2_90/Y vdd 6.82fF
C571 vdd DFFPOSX1_74/a_2_6# 5.17fF
C572 vdd DFFPOSX1_98/a_34_4# 2.60fF
C573 vdd OAI21X1_33/B 5.11fF
C574 vdd INVX2_49/Y 14.12fF
C575 DFFPOSX1_63/a_34_4# XOR2X1_81/A 2.07fF
C576 vdd XOR2X1_58/a_13_43# 2.11fF
C577 out_MuxData[9] out_MuxData[5] 3.39fF
C578 vdd XOR2X1_9/a_2_6# 2.07fF
C579 vdd XOR2X1_1/Y 11.64fF
C580 BUFX2_10/Y out_MemBData[13] 2.56fF
C581 XNOR2X1_45/A XNOR2X1_45/Y 2.02fF
C582 AOI22X1_99/Y vdd 11.42fF
C583 vdd XOR2X1_51/a_13_43# 2.11fF
C584 in_run vdd 9.21fF
C585 OR2X1_2/a_2_54# vdd 2.19fF
C586 XOR2X1_25/a_13_43# vdd 2.11fF
C587 DFFPOSX1_58/a_34_4# vdd 2.60fF
C588 vdd AND2X2_5/A 2.89fF
C589 vdd DFFPOSX1_0/a_34_4# 2.60fF
C590 vdd HAX1_4/a_2_74# 3.67fF
C591 vdd XOR2X1_16/a_13_43# 2.11fF
C592 vdd AOI22X1_0/a_2_54# 2.85fF
C593 vdd NAND3X1_34/Y 6.20fF
C594 vdd DFFPOSX1_8/a_22_6# 2.55fF
C595 INVX2_62/Y INVX2_106/Y 2.28fF
C596 gnd INVX2_94/Y 18.28fF
C597 INVX2_41/Y DFFPOSX1_20/a_22_6# 2.12fF
C598 XNOR2X1_30/a_12_41# AND2X2_38/Y 2.09fF
C599 OR2X2_0/A BUFX2_5/Y 2.41fF
C600 vdd XOR2X1_42/a_13_43# 2.11fF
C601 NAND2X1_6/Y vdd 5.75fF
C602 AOI22X1_13/a_2_54# vdd 2.85fF
C603 DFFPOSX1_5/a_2_6# vdd 5.17fF
C604 INVX2_93/A vdd 10.76fF
C605 DFFPOSX1_38/a_34_4# vdd 2.60fF
C606 gnd BUFX2_5/Y 29.96fF
C607 vdd INVX2_122/A 4.85fF
C608 vdd DFFPOSX1_37/a_2_6# 5.17fF
C609 vdd HAX1_13/B 7.21fF
C610 BUFX2_9/Y DFFPOSX1_28/a_22_6# 2.41fF
C611 vdd AOI22X1_52/a_2_54# 2.85fF
C612 vdd DFFPOSX1_4/a_2_6# 5.17fF
C613 vdd XOR2X1_28/a_2_6# 2.07fF
C614 vdd NAND3X1_14/A 2.85fF
C615 INVX2_5/A XNOR2X1_9/A 2.13fF
C616 XOR2X1_53/a_13_43# XOR2X1_17/B 3.65fF
C617 out_MuxData[15] out_MuxData[5] 2.13fF
C618 XOR2X1_2/a_13_43# vdd 2.11fF
C619 INVX2_86/A INVX2_67/A 2.84fF
C620 XNOR2X1_41/Y NAND2X1_28/Y 2.25fF
C621 XOR2X1_71/Y XNOR2X1_49/a_12_41# 2.64fF
C622 vdd DFFPOSX1_79/a_2_6# 5.17fF
C623 vdd INVX2_130/A 5.96fF
C624 vdd NAND3X1_3/Y 5.91fF
C625 con_count[3] gnd 6.25fF
C626 vdd OAI21X1_73/C 5.75fF
C627 AND2X2_36/B gnd 3.77fF
C628 NOR2X1_10/B vdd 3.96fF
C629 vdd INVX2_81/Y 2.62fF
C630 INVX2_86/A XOR2X1_55/B 3.00fF
C631 INVX2_56/A gnd 2.63fF
C632 out_MuxData[12] out_MuxData[10] 2.29fF
C633 INVX2_7/A INVX2_11/A 2.13fF
C634 AOI22X1_18/C gnd 2.33fF
C635 vdd OAI21X1_76/Y 2.93fF
C636 vdd DFFPOSX1_8/a_2_6# 5.17fF
C637 out_MemBData[0] INVX2_71/A 2.10fF
C638 vdd XNOR2X1_25/a_2_6# 2.29fF
C639 gnd out_MuxData[10] 11.78fF
C640 NAND3X1_25/B XOR2X1_69/B 2.42fF
C641 vdd XNOR2X1_24/a_2_6# 2.29fF
C642 vdd DFFPOSX1_6/a_2_6# 5.17fF
C643 vdd BUFX2_3/Y 9.29fF
C644 out_MuxData[4] out_MuxData[10] 2.91fF
C645 out_MuxData[4] XOR2X1_14/a_2_6# 2.57fF
C646 AND2X2_12/Y vdd 3.31fF
C647 vdd AOI22X1_10/a_2_54# 2.85fF
C648 INVX2_41/Y BUFX2_9/Y 2.20fF
C649 BUFX2_11/a_2_6# vdd 2.41fF
C650 vdd con_countWriteout[1] 20.20fF
C651 out_MuxData[12] gnd 13.99fF
C652 XOR2X1_13/a_13_43# AND2X2_8/A 2.25fF
C653 OAI21X1_40/A gnd 3.20fF
C654 vdd OAI21X1_84/Y 3.72fF
C655 vdd XOR2X1_38/a_2_6# 2.07fF
C656 vdd DFFPOSX1_85/a_22_6# 2.55fF
C657 vdd NAND3X1_4/B 7.00fF
C658 BUFX2_9/Y DFFPOSX1_14/a_22_6# 2.18fF
C659 vdd INVX2_30/Y 4.72fF
C660 AND2X2_19/Y gnd 13.21fF
C661 out_MuxData[4] gnd 8.73fF
C662 vdd XOR2X1_11/a_13_43# 2.11fF
C663 INVX2_41/Y DFFPOSX1_7/a_22_6# 3.34fF
C664 vdd XOR2X1_60/a_13_43# 2.11fF
C665 vdd DFFPOSX1_73/a_34_4# 2.60fF
C666 AOI22X1_7/a_2_54# vdd 2.85fF
C667 XNOR2X1_30/a_2_6# vdd 2.29fF
C668 INVX2_55/Y vdd 6.49fF
C669 NAND3X1_16/B AND2X2_16/Y 3.39fF
C670 vdd INVX2_3/Y 5.53fF
C671 vdd OAI21X1_80/C 3.88fF
C672 vdd XOR2X1_34/a_2_6# 2.07fF
C673 vdd XNOR2X1_4/a_2_6# 2.29fF
C674 vdd DFFPOSX1_31/a_22_6# 2.55fF
C675 INVX2_73/Y gnd 20.10fF
C676 vdd DFFPOSX1_96/a_2_6# 5.17fF
C677 vdd XOR2X1_7/Y 9.21fF
C678 OAI21X1_0/A out_MuxData[5] 2.09fF
C679 out_MuxData[3] out_MuxData[0] 2.60fF
C680 OAI21X1_68/B NOR2X1_28/B 2.04fF
C681 AND2X2_26/Y vdd 2.71fF
C682 INVX2_99/Y INVX2_84/Y 4.59fF
C683 vdd AOI22X1_10/C 2.68fF
C684 vdd XNOR2X1_2/a_2_6# 2.29fF
C685 vdd INVX2_39/A 19.89fF
C686 vdd AOI22X1_57/a_2_54# 2.85fF
C687 vdd DFFPOSX1_27/a_34_4# 2.60fF
C688 XOR2X1_76/Y AOI22X1_90/a_2_54# 2.03fF
C689 vdd INVX2_126/A 23.20fF
C690 vdd XOR2X1_88/B 4.27fF
C691 AND2X2_38/Y gnd 2.82fF
C692 vdd XOR2X1_40/A 6.07fF
C693 vdd DFFPOSX1_25/a_34_4# 2.60fF
C694 vdd NAND2X1_28/Y 10.10fF
C695 vdd AOI22X1_42/a_2_54# 2.85fF
C696 vdd INVX2_5/A 21.30fF
C697 vdd INVX2_52/A 18.15fF
C698 vdd DFFPOSX1_47/a_2_6# 5.17fF
C699 vdd AND2X2_24/Y 4.22fF
C700 NAND3X1_6/Y vdd 8.30fF
C701 AOI22X1_48/a_2_54# vdd 2.85fF
C702 INVX2_30/A vdd 5.06fF
C703 XOR2X1_66/a_13_43# vdd 2.11fF
C704 AOI22X1_55/Y vdd 3.18fF
C705 BUFX2_8/A out_MemBData[15] 2.48fF
C706 INVX2_93/Y gnd 2.96fF
C707 XOR2X1_81/A gnd 31.87fF
C708 vdd out_MuxData[2] 50.86fF
C709 vdd XNOR2X1_59/a_2_6# 2.29fF
C710 XOR2X1_67/a_13_43# vdd 2.11fF
C711 DFFPOSX1_5/a_2_6# con_countWriteout[4] 2.01fF
C712 out_state[2] vdd 11.57fF
C713 XNOR2X1_44/a_2_6# vdd 2.29fF
C714 out_MemBData[8] NOR2X1_48/Y 3.13fF
C715 NOR2X1_29/B vdd 2.97fF
C716 DFFPOSX1_55/a_2_6# INVX2_43/Y 2.35fF
C717 DFFPOSX1_70/a_34_4# vdd 2.60fF
C718 INVX2_5/A XOR2X1_46/a_2_6# 2.90fF
C719 OR2X1_0/a_2_54# vdd 2.19fF
C720 vdd DFFPOSX1_37/a_34_4# 2.60fF
C721 vdd OAI21X1_55/Y 2.51fF
C722 vdd XOR2X1_79/a_2_6# 2.07fF
C723 XOR2X1_23/A XNOR2X1_22/A 2.09fF
C724 vdd XOR2X1_91/a_13_43# 2.11fF
C725 vdd BUFX2_1/a_2_6# 2.41fF
C726 gnd XOR2X1_0/Y 2.26fF
C727 out_state[1] gnd 3.52fF
C728 INVX2_119/Y OR2X2_0/Y 3.17fF
C729 vdd OR2X2_0/Y 44.64fF
C730 DFFPOSX1_41/a_2_6# BUFX2_11/Y 2.82fF
C731 out_MemBData[3] vdd 17.80fF
C732 NAND2X1_4/A out_MuxData[15] 2.65fF
C733 vdd AND2X2_33/Y 3.43fF
C734 OAI21X1_2/A out_MuxData[14] 2.18fF
C735 vdd DFFPOSX1_45/a_2_6# 5.17fF
C736 vdd XOR2X1_50/a_13_43# 2.11fF
C737 vdd AOI22X1_91/a_2_54# 2.85fF
C738 out_MuxData[9] out_MuxData[0] 2.49fF
C739 vdd AOI22X1_79/a_2_54# 2.85fF
C740 out_MemBData[2] gnd 8.63fF
C741 AOI22X1_65/a_2_54# INVX2_94/Y 2.19fF
C742 vdd AOI22X1_48/D 2.12fF
C743 NOR2X1_9/Y AND2X2_17/A 2.01fF
C744 out_MuxData[1] vdd 52.26fF
C745 AOI21X1_2/B vdd 4.97fF
C746 INVX2_86/A gnd 2.15fF
C747 vdd INVX2_92/Y 46.00fF
C748 vdd out_win 8.14fF
C749 vdd DFFPOSX1_10/a_2_6# 5.17fF
C750 vdd AOI22X1_99/a_2_54# 2.85fF
C751 vdd DFFPOSX1_26/a_22_6# 2.55fF
C752 vdd out_MuxData[5] 87.89fF
C753 DFFPOSX1_31/a_34_4# NOR2X1_41/B 2.22fF
C754 XOR2X1_23/a_13_43# vdd 2.11fF
C755 DFFPOSX1_57/a_22_6# vdd 2.55fF
C756 BUFX2_10/Y gnd 22.54fF
C757 vdd DFFPOSX1_37/a_22_6# 2.55fF
C758 vdd AOI22X1_59/a_2_54# 2.85fF
C759 vdd BUFX2_1/Y 6.92fF
C760 BUFX2_10/Y out_MuxData[4] 4.26fF
C761 vdd XNOR2X1_45/Y 6.10fF
C762 vdd BUFX2_11/Y 81.72fF
C763 XNOR2X1_36/a_2_6# INVX2_28/Y 2.10fF
C764 vdd INVX2_25/Y 8.56fF
C765 NOR2X1_0/B XOR2X1_0/B 2.17fF
C766 vdd DFFPOSX1_100/a_22_6# 2.55fF
C767 vdd AOI22X1_44/a_2_54# 2.85fF
C768 vdd DFFPOSX1_11/a_2_6# 5.17fF
C769 vdd AOI22X1_37/a_2_54# 2.85fF
C770 INVX2_16/Y out_MuxData[10] 3.97fF
C771 XNOR2X1_32/a_2_6# XOR2X1_17/B 2.82fF
C772 AOI22X1_70/a_2_54# vdd 2.85fF
C773 DFFPOSX1_55/a_34_4# vdd 2.60fF
C774 vdd AND2X2_5/B 6.83fF
C775 vdd INVX2_53/A 11.99fF
C776 vdd OAI21X1_38/C 8.52fF
C777 INVX2_15/A INVX2_11/A 2.01fF
C778 vdd INVX2_43/Y 55.36fF
C779 vdd NAND2X1_10/Y 4.41fF
C780 vdd XOR2X1_38/a_13_43# 2.11fF
C781 vdd XOR2X1_18/a_13_43# 2.07fF
C782 INVX2_16/Y out_MuxData[12] 3.41fF
C783 vdd DFFPOSX1_19/a_22_6# 2.55fF
C784 con_count[1] con_count[0] 2.92fF
C785 INVX2_16/Y gnd 12.41fF
C786 vdd XOR2X1_57/a_13_43# 2.11fF
C787 INVX2_72/A vdd 4.20fF
C788 vdd INVX2_62/Y 37.33fF
C789 vdd DFFPOSX1_0/a_2_6# 5.17fF
C790 XOR2X1_64/B INVX2_28/Y 2.09fF
C791 XOR2X1_58/B gnd 2.24fF
C792 gnd AND2X2_13/Y 2.16fF
C793 AND2X2_20/Y gnd 2.35fF
C794 NOR2X1_49/B NOR2X1_49/Y 2.03fF
C795 DFFPOSX1_4/a_34_4# vdd 2.60fF
C796 BUFX2_9/Y DFFPOSX1_80/a_2_6# 2.05fF
C797 con_writeout gnd 5.58fF
C798 INVX2_97/Y vdd 3.28fF
C799 vdd NOR2X1_14/B 2.62fF
C800 NOR2X1_4/Y vdd 3.46fF
C801 vdd XOR2X1_23/A 2.48fF
C802 vdd DFFPOSX1_22/a_34_4# 2.60fF
C803 vdd DFFPOSX1_80/a_34_4# 2.60fF
C804 vdd XOR2X1_89/Y 7.91fF
C805 vdd AOI22X1_21/a_2_54# 2.85fF
C806 out_MuxData[10] out_MuxData[6] 4.73fF
C807 AND2X2_0/Y BUFX2_5/Y 2.37fF
C808 vdd AOI22X1_80/a_2_54# 2.85fF
C809 vdd out_MemBData[5] 14.59fF
C810 con_loseSig gnd 4.39fF
C811 vdd DFFPOSX1_54/a_2_6# 5.17fF
C812 vdd DFFPOSX1_83/a_34_4# 2.60fF
C813 INVX2_132/Y NOR2X1_47/B 2.44fF
C814 vdd AOI22X1_93/C 2.68fF
C815 vdd XNOR2X1_10/a_2_6# 2.29fF
C816 gnd out_MuxData[6] 4.47fF
C817 XOR2X1_7/a_13_43# vdd 2.11fF
C818 out_MuxData[4] out_MuxData[6] 4.67fF
C819 vdd XNOR2X1_38/a_2_6# 2.29fF
C820 vdd XNOR2X1_12/a_2_6# 2.29fF
C821 vdd NOR2X1_44/B 3.20fF
C822 XOR2X1_10/a_13_43# vdd 2.11fF
C823 XOR2X1_70/a_2_6# vdd 2.07fF
C824 AND2X2_36/A AND2X2_36/B 2.03fF
C825 vdd AOI22X1_34/a_2_54# 2.85fF
C826 vdd DFFPOSX1_17/a_2_6# 5.17fF
C827 vdd AOI21X1_3/Y 4.54fF
C828 INVX2_41/Y out_MemBData[3] 2.36fF
C829 INVX2_4/A vdd 3.63fF
C830 out_MuxData[7] out_MuxData[12] 3.08fF
C831 XOR2X1_10/a_2_6# out_MuxData[2] 3.52fF
C832 out_MuxData[7] gnd 13.38fF
C833 XNOR2X1_46/a_2_6# vdd 2.29fF
C834 vdd DFFPOSX1_15/a_34_4# 2.60fF
C835 vdd XNOR2X1_0/Y 11.43fF
C836 vdd DFFPOSX1_97/a_22_6# 2.55fF
C837 vdd XOR2X1_85/a_2_6# 2.07fF
C838 XOR2X1_60/a_13_43# INVX2_85/Y 2.64fF
C839 BUFX2_9/Y INVX2_11/A 2.10fF
C840 out_MemBData[5] INVX2_118/A 2.13fF
C841 vdd DFFPOSX1_44/a_34_4# 2.60fF
C842 vdd DFFPOSX1_43/a_34_4# 2.60fF
C843 vdd NOR2X1_5/Y 5.35fF
C844 gnd INVX2_71/Y 3.21fF
C845 XOR2X1_32/a_2_6# out_MuxData[5] 2.70fF
C846 NAND2X1_4/A vdd 2.89fF
C847 vdd DFFPOSX1_73/a_2_6# 5.17fF
C848 XOR2X1_13/a_13_43# vdd 2.11fF
C849 XOR2X1_29/a_13_43# vdd 2.11fF
C850 vdd XOR2X1_33/Y 3.20fF
C851 out_MuxData[12] NOR2X1_2/B 2.03fF
C852 vdd XOR2X1_62/B 2.21fF
C853 AND2X2_36/A gnd 4.73fF
C854 out_temp_addNum[0] BUFX2_2/Y 2.27fF
C855 vdd DFFPOSX1_87/a_22_6# 2.55fF
C856 INVX2_86/Y XOR2X1_47/a_13_43# 2.66fF
C857 con_count[8] gnd 6.51fF
C858 vdd XOR2X1_33/B 9.56fF
C859 vdd DFFPOSX1_52/a_34_4# 2.60fF
C860 vdd NAND2X1_3/A 5.43fF
C861 vdd XOR2X1_30/Y 4.50fF
C862 AOI22X1_9/a_2_54# vdd 2.85fF
C863 vdd NOR2X1_33/Y 3.61fF
C864 XOR2X1_41/a_2_6# INVX2_28/Y 2.80fF
C865 vdd XOR2X1_55/a_2_6# 2.07fF
C866 AND2X2_8/B vdd 11.52fF
C867 XOR2X1_66/Y vdd 2.91fF
C868 vdd XOR2X1_33/a_13_43# 2.11fF
C869 DFFPOSX1_41/a_22_6# BUFX2_11/Y 3.21fF
C870 vdd NOR2X1_45/A 4.47fF
C871 INVX2_72/Y AND2X2_35/a_2_6# 2.32fF
C872 vdd NOR2X1_15/B 6.16fF
C873 vdd DFFPOSX1_50/a_34_4# 2.60fF
C874 vdd INVX2_68/Y 7.36fF
C875 vdd OR2X1_1/a_2_54# 2.19fF
C876 vdd con_countWriteout[0] 11.05fF
C877 vdd DFFPOSX1_39/a_34_4# 2.60fF
C878 DFFPOSX1_60/a_2_6# vdd 5.13fF
C879 con_count[6] vdd 4.33fF
C880 OAI21X1_27/Y NAND2X1_9/Y 2.19fF
C881 vdd NOR2X1_49/B 2.24fF
C882 INVX2_126/Y con_count[4] 2.37fF
C883 vdd out_MuxData[0] 51.67fF
C884 vdd XNOR2X1_17/a_2_6# 2.29fF
C885 gnd NAND2X1_9/Y 4.70fF
C886 AOI22X1_71/a_2_54# vdd 2.85fF
C887 vdd AOI22X1_56/a_2_54# 2.85fF
C888 DFFPOSX1_70/a_2_6# vdd 5.17fF
C889 vdd con_count[2] 17.65fF
C890 vdd XOR2X1_76/Y 4.90fF
C891 vdd XNOR2X1_24/Y 7.23fF
C892 vdd XOR2X1_15/B 3.70fF
C893 out_MuxData[3] gnd 15.00fF
C894 vdd AND2X2_7/Y 3.03fF
C895 AND2X2_39/Y XOR2X1_69/B 2.92fF
C896 vdd NOR2X1_41/B 33.94fF
C897 vdd DFFPOSX1_13/a_2_6# 5.17fF
C898 XOR2X1_20/a_2_6# out_MuxData[4] 3.71fF
C899 vdd AND2X2_31/Y 3.90fF
C900 vdd NOR2X1_9/B 2.91fF
C901 vdd AOI22X1_15/a_2_54# 2.85fF
C902 XOR2X1_52/a_2_6# vdd 2.07fF
C903 out_temp_addNum[0] gnd 13.22fF
C904 vdd HAX1_3/YS 3.50fF
C905 vdd XOR2X1_88/a_2_6# 2.07fF
C906 vdd XOR2X1_0/a_13_43# 2.11fF
C907 vdd DFFPOSX1_51/a_34_4# 2.60fF
C908 DFFPOSX1_63/a_2_6# vdd 5.17fF
C909 XOR2X1_69/A gnd 4.57fF
C910 INVX2_93/A DFFPOSX1_67/a_34_4# 2.50fF
C911 vdd INVX2_59/A 8.14fF
C912 out_MuxData[8] INVX2_17/Y 2.42fF
C913 vdd DFFPOSX1_3/a_22_6# 2.55fF
C914 out_MuxData[11] out_MuxData[5] 2.34fF
C915 vdd DFFPOSX1_98/a_2_6# 5.17fF
C916 vdd NAND3X1_15/B 7.56fF
C917 gnd INVX2_106/Y 5.06fF
C918 OAI21X1_87/A gnd 2.47fF
C919 vdd DFFPOSX1_11/a_22_6# 2.55fF
C920 INVX2_11/Y con_countWriteout[5] 2.53fF
C921 vdd DFFPOSX1_75/a_34_4# 2.60fF
C922 vdd HAX1_9/B 5.52fF
C923 AOI22X1_96/Y gnd 5.19fF
C924 out_MemBData[1] vdd 19.75fF
C925 vdd con_count[0] 25.60fF
C926 vdd OAI21X1_57/C 5.24fF
C927 vdd XOR2X1_30/a_2_6# 2.07fF
C928 vdd DFFPOSX1_49/a_34_4# 2.60fF
C929 vdd DFFPOSX1_33/a_34_4# 2.60fF
C930 INVX2_16/Y out_MuxData[6] 2.43fF
C931 vdd DFFPOSX1_51/a_2_6# 5.17fF
C932 vdd NAND2X1_13/Y 10.83fF
C933 NOR2X1_44/A XNOR2X1_53/a_12_41# 2.55fF
C934 vdd out_MemBData[13] 6.31fF
C935 con_count[1] gnd 4.93fF
C936 out_MuxData[9] gnd 8.52fF
C937 vdd BUFX2_6/Y 6.52fF
C938 INVX2_61/Y INVX2_62/Y 3.67fF
C939 vdd DFFPOSX1_77/a_34_4# 2.60fF
C940 vdd INVX2_49/A 2.44fF
C941 vdd HAX1_2/a_2_74# 3.67fF
C942 vdd XOR2X1_54/a_13_43# 2.11fF
C943 vdd XOR2X1_36/B 6.12fF
C944 vdd XOR2X1_36/a_2_6# 2.07fF
C945 vdd XNOR2X1_60/a_2_6# 2.29fF
C946 OAI21X1_87/A INVX2_123/Y 2.04fF
C947 out_MuxData[2] out_MuxData[14] 2.49fF
C948 DFFPOSX1_58/a_2_6# vdd 5.17fF
C949 vdd NOR2X1_34/Y 12.18fF
C950 DFFPOSX1_40/a_34_4# out_MuxData[10] 2.27fF
C951 vdd in_clkb 27.07fF
C952 vdd NAND3X1_7/B 2.86fF
C953 vdd DFFPOSX1_91/a_22_6# 2.55fF
C954 INVX2_46/A gnd 2.03fF
C955 vdd XOR2X1_91/Y 4.62fF
C956 NAND3X1_15/Y OAI21X1_33/B 2.86fF
C957 OAI21X1_2/C XOR2X1_3/Y 4.99fF
C958 vdd INVX2_51/Y 4.13fF
C959 vdd OAI22X1_6/C 35.40fF
C960 vdd XOR2X1_29/a_2_6# 2.07fF
C961 vdd XOR2X1_44/a_13_43# 2.11fF
C962 gnd out_MuxData[15] 10.71fF
C963 vdd AOI22X1_99/B 3.04fF
C964 con_loadData con_readData 2.59fF
C965 out_MuxData[8] XOR2X1_65/Y 2.46fF
C966 out_MuxData[1] out_MuxData[14] 2.89fF
C967 vdd OAI21X1_45/C 3.88fF
C968 INVX2_67/A vdd 5.97fF
C969 DFFPOSX1_63/a_34_4# vdd 2.60fF
C970 XOR2X1_76/a_13_43# out_MuxData[2] 2.66fF
C971 vdd OAI21X1_73/Y 4.49fF
C972 vdd XOR2X1_41/A 2.08fF
C973 out_MuxData[7] out_MuxData[6] 2.45fF
C974 vdd AOI22X1_95/a_2_54# 2.85fF
C975 vdd XOR2X1_87/a_2_6# 2.07fF
C976 con_countWriteout[6] HAX1_1/a_2_74# 2.88fF
C977 INVX2_39/A XOR2X1_45/a_13_43# 3.65fF
C978 XOR2X1_1/B OAI21X1_2/A 2.33fF
C979 XOR2X1_23/a_13_43# out_MuxData[14] 2.58fF
C980 XOR2X1_51/a_13_43# INVX2_87/Y 3.65fF
C981 con_countWriteout[0] AOI22X1_29/a_2_54# 2.06fF
C982 DFFPOSX1_35/a_2_6# INVX2_43/Y 2.42fF
C983 XOR2X1_63/Y XNOR2X1_45/Y 3.05fF
C984 XOR2X1_70/a_13_43# vdd 2.11fF
C985 vdd XOR2X1_33/a_2_6# 2.07fF
C986 vdd AND2X2_41/A 7.26fF
C987 vdd DFFPOSX1_8/a_34_4# 2.60fF
C988 vdd XOR2X1_55/B 11.68fF
C989 vdd DFFPOSX1_92/a_34_4# 2.60fF
C990 vdd AOI22X1_87/C 2.68fF
C991 vdd AOI22X1_55/a_2_54# 2.85fF
C992 vdd XOR2X1_28/a_13_43# 2.11fF
C993 AOI21X1_6/B out_MuxData[10] 2.74fF
C994 AOI22X1_3/a_2_54# vdd 2.85fF
C995 INVX2_11/Y gnd 5.34fF
C996 vdd XOR2X1_51/Y 2.97fF
C997 XOR2X1_74/Y out_MuxData[0] 3.15fF
C998 XOR2X1_20/a_13_43# vdd 2.11fF
C999 XNOR2X1_21/a_2_6# vdd 2.29fF
C1000 OAI22X1_6/C XNOR2X1_54/a_2_6# 2.28fF
C1001 INVX2_60/Y vdd 4.88fF
C1002 OAI21X1_91/A gnd 2.00fF
C1003 NOR2X1_29/A gnd 2.21fF
C1004 vdd INVX2_72/Y 25.72fF
C1005 vdd con_countWriteout[5] 10.01fF
C1006 vdd DFFPOSX1_97/a_34_4# 2.60fF
C1007 vdd DFFPOSX1_17/a_22_6# 2.55fF
C1008 out_MuxData[1] XNOR2X1_22/a_12_41# 2.45fF
C1009 vdd NAND3X1_16/A 5.24fF
C1010 vdd INVX2_73/A 10.91fF
C1011 vdd DFFPOSX1_85/a_34_4# 2.60fF
C1012 vdd XOR2X1_8/a_2_6# 2.07fF
C1013 DFFPOSX1_36/a_2_6# vdd 5.17fF
C1014 XOR2X1_68/a_2_6# vdd 2.07fF
C1015 out_MemBData[12] vdd 23.93fF
C1016 OAI21X1_69/C vdd 2.78fF
C1017 INVX2_41/Y DFFPOSX1_3/a_22_6# 2.16fF
C1018 out_MuxData[1] XOR2X1_78/a_2_6# 2.22fF
C1019 vdd DFFPOSX1_19/a_34_4# 2.60fF
C1020 vdd AOI22X1_45/a_2_54# 2.85fF
C1021 XOR2X1_63/a_13_43# vdd 2.11fF
C1022 XNOR2X1_48/a_12_41# XOR2X1_77/Y 2.78fF
C1023 vdd DFFPOSX1_87/a_34_4# 2.60fF
C1024 vdd AOI22X1_17/a_2_54# 2.85fF
C1025 vdd AOI22X1_63/a_2_54# 2.85fF
C1026 vdd AOI22X1_61/B 9.68fF
C1027 vdd OAI22X1_11/Y 2.82fF
C1028 vdd XOR2X1_34/a_13_43# 2.11fF
C1029 vdd XOR2X1_26/Y 5.26fF
C1030 vdd AOI22X1_8/a_2_54# 2.85fF
C1031 con_restart OR2X2_0/Y 2.22fF
C1032 INVX2_34/Y gnd 2.56fF
C1033 vdd NOR2X1_42/B 4.18fF
C1034 AOI22X1_68/a_2_54# vdd 2.85fF
C1035 vdd AOI22X1_46/a_2_54# 2.85fF
C1036 vdd INVX2_6/A 2.59fF
C1037 DFFPOSX1_68/a_22_6# vdd 2.55fF
C1038 XOR2X1_43/a_13_43# vdd 2.11fF
C1039 vdd NAND3X1_1/B 4.14fF
C1040 vdd BUFX2_2/Y 27.47fF
C1041 INVX2_86/Y XOR2X1_57/a_13_43# 2.06fF
C1042 vdd AOI22X1_86/a_2_54# 2.85fF
C1043 vdd DFFPOSX1_25/a_2_6# 5.17fF
C1044 vdd DFFPOSX1_94/a_22_6# 2.55fF
C1045 vdd XOR2X1_16/a_2_6# 2.07fF
C1046 vdd XOR2X1_27/a_2_6# 2.07fF
C1047 vdd INVX2_10/Y 4.76fF
C1048 OAI21X1_75/Y BUFX2_11/Y 2.01fF
C1049 vdd INVX2_94/Y 15.08fF
C1050 BUFX2_4/Y gnd 13.79fF
C1051 XOR2X1_2/Y gnd 4.10fF
C1052 XOR2X1_69/A OAI21X1_89/A 2.13fF
C1053 vdd XOR2X1_2/a_2_6# 2.07fF
C1054 vdd AND2X2_28/A 8.31fF
C1055 out_MuxData[11] out_MuxData[0] 4.39fF
C1056 vdd BUFX2_5/Y 64.33fF
C1057 AND2X2_11/a_2_6# AND2X2_6/B 2.51fF
C1058 out_MuxData[1] XOR2X1_17/B 2.23fF
C1059 XOR2X1_62/a_2_6# vdd 2.07fF
C1060 vdd AOI22X1_59/C 2.68fF
C1061 con_count[8] INVX2_70/A 2.64fF
C1062 vdd DFFPOSX1_2/a_34_4# 2.60fF
C1063 INVX2_88/Y INVX2_43/Y 2.61fF
C1064 vdd con_count[3] 16.26fF
C1065 NAND3X1_3/C XOR2X1_26/a_2_6# 2.17fF
C1066 vdd DFFPOSX1_47/a_34_4# 2.60fF
C1067 XOR2X1_40/A XOR2X1_40/a_2_6# 2.65fF
C1068 XOR2X1_48/B out_MuxData[3] 2.58fF
C1069 vdd AND2X2_36/B 8.36fF
C1070 vdd DFFPOSX1_17/a_34_4# 2.60fF
C1071 INVX2_21/A vdd 7.84fF
C1072 DFFPOSX1_57/a_2_6# vdd 5.17fF
C1073 XOR2X1_73/a_13_43# XOR2X1_81/A 2.64fF
C1074 vdd HAX1_5/a_2_74# 3.67fF
C1075 HAX1_3/B vdd 4.44fF
C1076 vdd INVX2_56/A 5.01fF
C1077 vdd XOR2X1_77/a_2_6# 2.07fF
C1078 AOI22X1_18/C vdd 2.68fF
C1079 XNOR2X1_39/a_2_6# vdd 2.29fF
C1080 OAI21X1_38/C con_restart 2.79fF
C1081 vdd INVX2_80/Y 3.36fF
C1082 vdd NOR2X1_46/B 46.83fF
C1083 vdd XOR2X1_65/a_2_6# 2.07fF
C1084 vdd out_MuxData[10] 58.99fF
C1085 vdd XOR2X1_88/a_13_43# 2.11fF
C1086 vdd INVX2_71/A 4.40fF
C1087 vdd INVX2_135/Y 3.44fF
C1088 vdd DFFPOSX1_33/a_2_6# 5.17fF
C1089 vdd XOR2X1_84/a_2_6# 2.07fF
C1090 XNOR2X1_8/a_2_6# XOR2X1_0/Y 2.96fF
C1091 vdd AND2X2_39/A 4.91fF
C1092 vdd XOR2X1_14/a_2_6# 2.07fF
C1093 vdd XOR2X1_22/a_2_6# 2.07fF
C1094 XNOR2X1_59/a_2_6# OAI21X1_90/Y 2.10fF
C1095 BUFX2_2/a_2_6# vdd 2.41fF
C1096 vdd OAI21X1_27/Y 2.22fF
C1097 out_MuxData[12] vdd 77.53fF
C1098 out_MemBData[0] vdd 9.57fF
C1099 vdd OAI21X1_40/A 5.06fF
C1100 vdd gnd 28.70fF
C1101 XNOR2X1_46/a_2_6# INVX2_86/Y 2.10fF
C1102 vdd DFFPOSX1_26/a_34_4# 2.60fF
C1103 vdd AND2X2_19/Y 44.40fF
C1104 vdd out_MuxData[4] 85.78fF
C1105 DFFPOSX1_57/a_34_4# vdd 2.60fF
C1106 vdd DFFPOSX1_75/a_2_6# 5.17fF
C1107 vdd DFFPOSX1_34/a_22_6# 2.55fF
C1108 vdd XOR2X1_80/a_2_6# 2.07fF
C1109 vdd INVX2_9/Y 2.25fF
C1110 vdd DFFPOSX1_95/a_22_6# 2.55fF
C1111 vdd INVX2_73/Y 10.47fF
C1112 vdd DFFPOSX1_84/a_22_6# 2.55fF
C1113 vdd AOI22X1_50/a_2_54# 2.85fF
C1114 vdd DFFPOSX1_16/a_22_6# 2.55fF
C1115 NAND2X1_5/Y vdd 10.31fF
C1116 DFFPOSX1_14/a_34_4# vdd 2.60fF
C1117 XOR2X1_73/a_2_6# vdd 2.07fF
C1118 vdd AOI22X1_6/a_2_54# 2.85fF
C1119 INVX2_41/Y DFFPOSX1_17/a_22_6# 2.05fF
C1120 vdd AND2X2_38/Y 24.63fF
C1121 vdd DFFPOSX1_62/a_34_4# 2.60fF
C1122 vdd OAI21X1_69/Y 2.37fF
C1123 vdd DFFPOSX1_22/a_2_6# 5.17fF
C1124 vdd INVX2_123/Y 7.11fF
C1125 NOR2X1_16/B gnd 2.30fF
C1126 AND2X2_7/Y con_countWriteout[2] 2.74fF
C1127 BUFX2_8/A INVX2_60/Y 2.30fF
C1128 OAI21X1_71/Y OAI21X1_71/C 2.05fF
C1129 INVX2_16/Y XOR2X1_19/a_2_6# 2.54fF
C1130 vdd XOR2X1_45/a_2_6# 2.07fF
C1131 vdd XOR2X1_57/A 3.99fF
C1132 AOI22X1_75/a_2_54# vdd 2.85fF
C1133 vdd AND2X2_17/A 5.59fF
C1134 AOI22X1_41/Y out_MuxData[13] 2.47fF
C1135 vdd INVX2_93/Y 37.78fF
C1136 vdd AOI22X1_35/a_2_54# 2.85fF
C1137 vdd XNOR2X1_57/a_2_6# 2.29fF
C1138 INVX2_10/A gnd 4.48fF
C1139 vdd XOR2X1_81/A 39.31fF
C1140 AOI22X1_34/a_2_54# INVX2_59/Y 2.03fF
C1141 vdd XOR2X1_14/a_13_43# 2.11fF
C1142 vdd XOR2X1_86/a_2_6# 2.07fF
C1143 out_MuxData[1] out_MuxData[8] 2.39fF
C1144 XNOR2X1_3/a_2_6# vdd 2.29fF
C1145 AOI22X1_78/a_2_54# vdd 2.85fF
C1146 vdd DFFPOSX1_62/a_22_6# 2.55fF
C1147 vdd AOI22X1_39/a_2_54# 2.85fF
C1148 vdd XOR2X1_0/Y 13.09fF
C1149 vdd out_state[1] 19.74fF
C1150 BUFX2_10/Y DFFPOSX1_74/a_22_6# 2.21fF
C1151 BUFX2_3/Y AOI22X1_38/A 2.03fF
C1152 INVX2_41/Y BUFX2_5/Y 2.56fF
C1153 vdd XOR2X1_61/a_2_6# 2.07fF
C1154 INVX2_84/Y out_MuxData[5] 4.58fF
C1155 vdd out_MemBData[2] 5.43fF
C1156 vdd DFFPOSX1_24/a_22_6# 2.55fF
C1157 vdd DFFPOSX1_82/a_34_4# 2.60fF
C1158 vdd INVX2_12/Y 2.85fF
C1159 vdd XOR2X1_18/B 3.17fF
C1160 AND2X2_21/A AOI22X1_55/Y 2.25fF
C1161 XNOR2X1_22/A out_MuxData[6] 2.04fF
C1162 NAND3X1_8/C XOR2X1_40/a_13_43# 2.63fF
C1163 INVX2_84/Y BUFX2_11/Y 2.98fF
C1164 AOI22X1_67/a_2_54# vdd 2.85fF
C1165 DFFPOSX1_35/a_22_6# INVX2_43/Y 2.09fF
C1166 INVX2_86/A vdd 33.06fF
C1167 DFFPOSX1_22/a_22_6# BUFX2_11/Y 2.44fF
C1168 vdd XOR2X1_23/a_2_6# 2.07fF
C1169 vdd DFFPOSX1_92/a_2_6# 5.17fF
C1170 INVX2_61/Y DFFPOSX1_97/a_34_4# 2.60fF
C1171 vdd AOI22X1_60/a_2_54# 2.85fF
C1172 vdd DFFPOSX1_80/a_22_6# 2.55fF
C1173 vdd INVX2_133/A 2.44fF
C1174 vdd XOR2X1_90/Y 4.61fF
C1175 OAI22X1_6/Y vdd 3.05fF
C1176 BUFX2_10/Y vdd 68.15fF
C1177 vdd DFFPOSX1_79/a_22_6# 2.55fF
C1178 BUFX2_9/a_2_6# vdd 2.41fF
C1179 con_countWriteout[4] gnd 3.25fF
C1180 NAND3X1_16/B out_MuxData[2] 2.97fF
C1181 vdd DFFPOSX1_97/a_2_6# 5.17fF
C1182 vdd NAND3X1_3/C 7.24fF
C1183 vdd XNOR2X1_22/a_2_6# 2.29fF
C1184 vdd DFFPOSX1_85/a_2_6# 5.17fF
C1185 vdd DFFPOSX1_43/a_2_6# 5.17fF
C1186 XOR2X1_63/a_2_6# vdd 2.07fF
C1187 XOR2X1_68/a_13_43# vdd 2.11fF
C1188 XOR2X1_25/a_2_6# vdd 2.07fF
C1189 AOI21X1_4/C vdd 4.31fF
C1190 vdd DFFPOSX1_78/a_2_6# 5.17fF
C1191 INVX2_41/Y gnd 14.75fF
C1192 DFFPOSX1_65/a_34_4# vdd 2.60fF
C1193 XNOR2X1_11/a_2_6# vdd 2.29fF
C1194 HAX1_3/B HAX1_3/a_41_74# 2.27fF
C1195 AOI22X1_88/C gnd 2.34fF
C1196 vdd AOI22X1_88/a_2_54# 2.85fF
C1197 DFFPOSX1_68/a_22_6# INVX2_61/Y 2.09fF
C1198 vdd XOR2X1_64/a_2_6# 2.07fF
C1199 out_state[0] gnd 3.87fF
C1200 vdd NAND3X1_17/B 9.46fF
C1201 vdd NOR2X1_21/Y 15.75fF
C1202 XOR2X1_76/a_2_6# out_MuxData[4] 4.38fF
C1203 INVX2_28/Y AND2X2_18/Y 3.39fF
C1204 INVX2_99/Y OAI22X1_9/Y 2.19fF
C1205 INVX2_99/A gnd 2.31fF
C1206 vdd XOR2X1_30/a_13_43# 2.11fF
C1207 vdd XOR2X1_38/Y 5.24fF
C1208 out_MuxData[11] NOR2X1_42/B 2.90fF
C1209 vdd NAND3X1_29/Y 7.01fF
C1210 INVX2_16/Y vdd 49.25fF
C1211 XNOR2X1_15/a_2_6# vdd 2.29fF
C1212 AOI22X1_68/C vdd 2.68fF
C1213 vdd AOI22X1_82/a_2_54# 2.85fF
C1214 INVX2_59/A INVX2_25/A 2.55fF
C1215 DFFPOSX1_68/a_34_4# vdd 2.60fF
C1216 vdd OAI22X1_17/Y 3.42fF
C1217 vdd XOR2X1_84/B 4.57fF
C1218 vdd XOR2X1_58/B 6.89fF
C1219 vdd AOI22X1_65/a_2_54# 2.85fF
C1220 vdd AND2X2_13/Y 14.19fF
C1221 vdd INVX2_129/Y 7.56fF
C1222 vdd AND2X2_20/Y 7.65fF
C1223 vdd DFFPOSX1_50/a_2_6# 5.17fF
C1224 vdd DFFPOSX1_42/a_22_6# 2.55fF
C1225 XOR2X1_70/Y XOR2X1_69/B 2.24fF
C1226 XNOR2X1_41/Y OAI21X1_58/Y 2.39fF
C1227 vdd AND2X2_13/B 2.54fF
C1228 AOI22X1_80/B vdd 6.85fF
C1229 OAI21X1_89/A vdd 9.75fF
C1230 AOI22X1_38/A OR2X2_0/Y 2.03fF
C1231 vdd XOR2X1_75/Y 2.30fF
C1232 vdd DFFPOSX1_39/a_2_6# 5.17fF
C1233 con_writeout vdd 28.28fF
C1234 INVX2_96/Y vdd 5.10fF
C1235 vdd INVX2_37/Y 6.82fF
C1236 INVX2_133/Y gnd 2.21fF
C1237 vdd AOI22X1_38/a_2_54# 2.85fF
C1238 vdd INVX2_135/A 4.00fF
C1239 vdd XOR2X1_1/a_2_6# 2.07fF
C1240 XOR2X1_12/a_2_6# vdd 2.07fF
C1241 BUFX2_9/Y DFFPOSX1_16/a_34_4# 2.70fF
C1242 XOR2X1_27/Y vdd 2.28fF
C1243 XOR2X1_46/a_2_6# AND2X2_13/Y 2.02fF
C1244 vdd HAX1_1/YS 3.00fF
C1245 vdd NOR2X1_15/A 8.12fF
C1246 vdd con_loseSig 15.11fF
C1247 vdd XOR2X1_65/A 2.87fF
C1248 vdd XOR2X1_83/a_2_6# 2.07fF
C1249 vdd AOI22X1_41/a_2_54# 2.85fF
C1250 vdd out_MuxData[6] 54.56fF
C1251 BUFX2_8/A INVX2_93/Y 2.83fF
C1252 DFFPOSX1_56/a_34_4# vdd 2.60fF
C1253 INVX2_66/A vdd 3.19fF
C1254 XOR2X1_52/a_13_43# vdd 2.11fF
C1255 vdd NOR2X1_48/B 29.81fF
C1256 vdd AOI22X1_96/a_2_54# 2.85fF
C1257 vdd HAX1_3/a_2_74# 3.67fF
C1258 INVX2_61/Y gnd 19.69fF
C1259 vdd XOR2X1_84/a_13_43# 2.11fF
C1260 INVX2_44/A gnd 16.78fF
C1261 vdd XOR2X1_56/a_2_6# 2.07fF
C1262 INVX2_85/Y gnd 2.12fF
C1263 out_MuxData[12] out_MuxData[11] 2.05fF
C1264 out_MuxData[11] NOR2X1_28/A 2.60fF
C1265 out_MuxData[11] gnd 14.10fF
C1266 out_MuxData[7] vdd 73.06fF
C1267 NOR2X1_22/Y gnd 2.77fF
C1268 vdd OAI21X1_4/A 6.56fF
C1269 in_clkb INVX2_59/Y 4.35fF
C1270 vdd XOR2X1_48/a_2_6# 2.07fF
C1271 gnd AND2X2_21/Y 10.75fF
C1272 vdd INVX2_71/Y 42.09fF
C1273 vdd OAI21X1_58/Y 4.37fF
C1274 vdd DFFPOSX1_11/a_34_4# 2.60fF
C1275 NOR2X1_28/B AOI22X1_57/a_2_54# 2.13fF
C1276 AOI22X1_64/a_2_54# vdd 2.85fF
C1277 vdd AND2X2_0/Y 2.95fF
C1278 XNOR2X1_16/a_2_6# XOR2X1_81/A 2.94fF
C1279 vdd AOI22X1_19/C 2.68fF
C1280 AND2X2_36/A vdd 14.99fF
C1281 vdd OAI21X1_44/C 8.46fF
C1282 vdd con_count[8] 10.77fF
C1283 vdd HAX1_6/a_2_74# 3.67fF
C1284 vdd XOR2X1_78/Y 5.44fF
C1285 vdd DFFPOSX1_95/a_34_4# 2.60fF
C1286 vdd DFFPOSX1_49/a_2_6# 5.17fF
C1287 XOR2X1_19/a_13_43# INVX2_17/Y 2.07fF
C1288 BUFX2_9/Y DFFPOSX1_92/a_22_6# 2.22fF
C1289 vdd DFFPOSX1_100/a_34_4# 2.60fF
C1290 vdd DFFPOSX1_30/a_22_6# 2.55fF
C1291 vdd DFFPOSX1_84/a_34_4# 2.60fF
C1292 con_countWriteout[7] DFFPOSX1_1/a_2_6# 2.05fF
C1293 BUFX2_4/a_2_6# vdd 2.41fF
C1294 vdd DFFPOSX1_19/a_2_6# 5.17fF
C1295 XOR2X1_35/a_2_6# vdd 2.07fF
C1296 vdd AOI22X1_60/C 2.68fF
C1297 vdd DFFPOSX1_50/a_22_6# 2.55fF
C1298 vdd NOR2X1_13/Y 5.55fF
C1299 NAND2X1_8/Y out_MuxData[4] 2.13fF
C1300 vdd out_temp_addNum[2] 3.89fF
C1301 INVX2_51/A gnd 2.56fF
C1302 XOR2X1_60/a_2_6# XOR2X1_81/A 2.44fF
C1303 vdd XOR2X1_6/a_2_6# 2.07fF
C1304 vdd XOR2X1_53/a_2_6# 2.07fF
C1305 BUFX2_10/Y INVX2_110/A 3.01fF
C1306 vdd INVX2_53/Y 2.48fF
C1307 XOR2X1_66/Y XNOR2X1_40/a_12_41# 2.75fF
C1308 HAX1_7/B vdd 6.83fF
C1309 INVX2_50/Y INVX2_17/Y 2.89fF
C1310 vdd XNOR2X1_50/a_2_6# 2.29fF
C1311 vdd XNOR2X1_52/a_2_6# 2.29fF
C1312 OAI21X1_67/Y vdd 3.06fF
C1313 vdd INVX2_48/Y 12.90fF
C1314 vdd DFFPOSX1_10/a_34_4# 2.60fF
C1315 vdd INVX2_70/A 13.33fF
C1316 vdd INVX2_65/A 4.85fF
C1317 AOI22X1_35/a_2_54# AND2X2_21/Y 2.03fF
C1318 vdd HAX1_12/B 6.17fF
C1319 vdd NAND2X1_9/Y 3.78fF
C1320 vdd DFFPOSX1_91/a_34_4# 2.60fF
C1321 vdd out_MemBData[6] 13.99fF
C1322 DFFPOSX1_53/a_34_4# out_MuxData[10] 2.06fF
C1323 INVX2_12/A vdd 4.09fF
C1324 vdd XOR2X1_15/a_13_43# 2.11fF
C1325 XOR2X1_74/B vdd 2.88fF
C1326 vdd AOI22X1_90/a_2_54# 2.85fF
C1327 AOI22X1_13/a_2_54# XOR2X1_19/Y 2.30fF
C1328 gnd con_countWriteout[2] 2.20fF
C1329 HAX1_13/a_41_74# INVX2_72/Y 2.10fF
C1330 vdd XOR2X1_20/a_2_6# 2.07fF
C1331 vdd out_MuxData[3] 22.45fF
C1332 BUFX2_9/Y DFFPOSX1_28/a_2_6# 2.17fF
C1333 out_MuxData[14] out_MuxData[10] 2.57fF
C1334 AND2X2_7/a_2_6# AND2X2_6/B 2.31fF
C1335 DFFPOSX1_36/a_34_4# vdd 2.60fF
C1336 NOR2X1_42/A vdd 6.63fF
C1337 INVX2_67/Y vdd 5.64fF
C1338 vdd INVX2_109/A 2.44fF
C1339 INVX2_99/Y OAI22X1_14/Y 2.16fF
C1340 vdd HAX1_5/YS 2.91fF
C1341 vdd out_temp_addNum[0] 3.97fF
C1342 vdd XOR2X1_11/a_2_6# 2.07fF
C1343 vdd AND2X2_8/A 3.25fF
C1344 gnd out_MuxData[14] 20.93fF
C1345 vdd DFFPOSX1_83/a_2_6# 5.17fF
C1346 vdd DFFPOSX1_82/a_2_6# 5.17fF
C1347 out_MuxData[4] out_MuxData[14] 2.18fF
C1348 OAI21X1_28/A vdd 8.13fF
C1349 XOR2X1_69/A vdd 25.87fF
C1350 HAX1_12/a_41_74# INVX2_126/A 2.02fF
C1351 NOR2X1_30/Y vdd 20.94fF
C1352 HAX1_2/B vdd 7.49fF
C1353 DFFPOSX1_69/a_22_6# vdd 2.55fF
C1354 AND2X2_29/Y vdd 3.42fF
C1355 vdd INVX2_19/A 11.51fF
C1356 vdd INVX2_106/Y 25.36fF
C1357 vdd DFFPOSX1_99/a_22_6# 2.55fF
C1358 vdd OAI21X1_87/A 5.70fF
C1359 INVX2_86/Y gnd 9.09fF
C1360 INVX2_15/Y out_MemBData[3] 3.17fF
C1361 vdd DFFPOSX1_79/a_34_4# 2.60fF
C1362 vdd AOI22X1_96/Y 8.89fF
C1363 vdd XOR2X1_49/Y 11.58fF
C1364 vdd DFFPOSX1_54/a_22_6# 2.55fF
C1365 INVX2_31/Y vdd 6.85fF
C1366 vdd INVX2_6/Y 5.73fF
C1367 vdd XOR2X1_11/Y 3.29fF
C1368 vdd XOR2X1_27/a_13_43# 2.11fF
C1369 vdd XOR2X1_17/a_13_43# 2.11fF
C1370 vdd DFFPOSX1_30/a_2_6# 5.17fF
C1371 vdd DFFPOSX1_46/a_22_6# 2.55fF
C1372 vdd OAI22X1_3/C 8.86fF
C1373 XOR2X1_37/a_2_6# out_MuxData[5] 2.65fF
C1374 BUFX2_3/a_2_6# vdd 2.41fF
C1375 vdd AND2X2_30/Y 4.58fF
C1376 INVX2_50/Y XOR2X1_65/Y 2.79fF
C1377 vdd DFFPOSX1_59/a_34_4# 2.60fF
C1378 vdd OAI22X1_16/Y 5.11fF
C1379 con_count[1] vdd 10.78fF
C1380 vdd XOR2X1_52/Y 3.85fF
C1381 DFFPOSX1_65/a_2_6# vdd 5.17fF
C1382 OAI21X1_79/C AND2X2_38/Y 3.20fF
C1383 vdd out_MuxData[9] 48.68fF
C1384 INVX2_11/A gnd 2.54fF
C1385 vdd AOI22X1_51/a_2_54# 2.85fF
C1386 vdd DFFPOSX1_31/a_34_4# 2.60fF
C1387 vdd NAND3X1_5/Y 3.61fF
C1388 INVX2_44/A AND2X2_20/Y 2.82fF
C1389 vdd AND2X2_38/B 2.03fF
C1390 AOI22X1_9/C vdd 2.68fF
C1391 DFFPOSX1_68/a_2_6# vdd 5.17fF
C1392 DFFPOSX1_23/a_2_6# vdd 5.17fF
C1393 con_writeout INVX2_61/Y 3.08fF
C1394 vdd XNOR2X1_49/a_2_6# 2.29fF
C1395 vdd AOI22X1_16/a_2_54# 2.85fF
C1396 vdd DFFPOSX1_94/a_34_4# 2.60fF
C1397 INVX2_126/Y INVX2_126/A 4.08fF
C1398 vdd XOR2X1_5/a_13_43# 2.11fF
C1399 vdd INVX2_134/A 2.44fF
C1400 INVX2_25/A gnd 3.36fF
C1401 vdd INVX2_46/A 14.76fF
C1402 vdd DFFPOSX1_25/a_22_6# 2.55fF
C1403 vdd XOR2X1_37/a_13_43# 2.11fF
C1404 NOR2X1_27/Y AOI21X1_6/B 3.41fF
C1405 XOR2X1_6/a_13_43# out_MuxData[6] 2.64fF
C1406 XNOR2X1_29/a_2_6# vdd 2.29fF
C1407 vdd DFFPOSX1_72/a_2_6# 5.13fF
C1408 vdd DFFPOSX1_89/a_22_6# 2.55fF
C1409 vdd XOR2X1_87/A 9.18fF
C1410 INVX2_57/A vdd 5.65fF
C1411 DFFPOSX1_40/a_34_4# vdd 2.60fF
C1412 DFFPOSX1_72/a_34_4# INVX2_126/A 2.37fF
C1413 vdd XNOR2X1_6/B 4.00fF
C1414 vdd XOR2X1_39/Y 2.39fF
C1415 vdd DFFPOSX1_3/a_34_4# 2.60fF
C1416 gnd con_restart 27.01fF
C1417 XOR2X1_4/Y out_MuxData[10] 2.49fF
C1418 vdd XOR2X1_21/a_2_6# 2.07fF
C1419 vdd XOR2X1_26/a_2_6# 2.07fF
C1420 XOR2X1_17/B out_MuxData[10] 2.04fF
C1421 vdd DFFPOSX1_53/a_22_6# 2.55fF
C1422 vdd out_MuxData[15] 47.67fF
C1423 vdd XOR2X1_32/a_13_43# 2.11fF
C1424 AND2X2_19/Y con_restart 3.10fF
C1425 INVX2_43/Y AND2X2_35/Y 2.88fF
C1426 INVX2_27/A vdd 5.09fF
C1427 DFFPOSX1_55/a_22_6# INVX2_43/Y 2.84fF
C1428 OAI21X1_68/A vdd 8.24fF
C1429 vdd INVX2_65/Y 6.10fF
C1430 XOR2X1_17/B gnd 11.36fF
C1431 XOR2X1_87/A AND2X2_37/a_2_6# 2.15fF
C1432 vdd DFFPOSX1_32/a_22_6# 2.55fF
C1433 vdd HAX1_6/YS 3.22fF
C1434 XOR2X1_8/a_13_43# out_MuxData[2] 2.47fF
C1435 OAI21X1_69/C out_MemBData[9] 2.26fF
C1436 NAND3X1_27/B vdd 4.47fF
C1437 DFFPOSX1_40/a_22_6# vdd 2.55fF
C1438 vdd DFFPOSX1_34/a_2_6# 5.17fF
C1439 XNOR2X1_8/A XNOR2X1_8/Y 2.09fF
C1440 vdd XOR2X1_77/a_13_43# 2.11fF
C1441 vdd NOR2X1_39/Y 10.79fF
C1442 vdd OAI21X1_89/B 11.87fF
C1443 vdd OAI21X1_81/Y 6.59fF
C1444 vdd XOR2X1_88/Y 4.90fF
C1445 vdd NOR2X1_8/A 4.22fF
C1446 OAI21X1_52/C INVX2_43/Y 2.10fF
C1447 vdd INVX2_125/Y 2.69fF
C1448 AOI22X1_67/a_2_54# con_count[7] 2.53fF
C1449 DFFPOSX1_2/a_22_6# BUFX2_5/Y 2.18fF
C1450 out_MuxData[7] out_MuxData[11] 2.17fF
C1451 OAI21X1_6/B XOR2X1_24/A 2.03fF
C1452 INVX2_11/Y vdd 24.25fF
C1453 INVX2_32/Y out_state[2] 2.11fF
C1454 vdd HAX1_9/YS 3.27fF
C1455 vdd OAI21X1_91/A 10.45fF
C1456 vdd XOR2X1_19/a_2_6# 2.07fF
C1457 INVX2_26/A gnd 2.72fF
C1458 vdd AOI22X1_93/a_2_54# 2.85fF
C1459 NAND2X1_8/Y out_MuxData[6] 2.79fF
C1460 vdd XOR2X1_39/a_13_43# 2.11fF
C1461 vdd XNOR2X1_22/A 4.04fF
C1462 vdd DFFPOSX1_47/a_22_6# 2.55fF
C1463 vdd DFFPOSX1_26/a_2_6# 5.17fF
C1464 XOR2X1_45/Y INVX2_46/A 2.46fF
C1465 vdd AOI21X1_6/B 4.64fF
C1466 vdd DFFPOSX1_3/a_2_6# 5.17fF
C1467 AOI22X1_3/C vdd 2.68fF
C1468 vdd DFFPOSX1_34/a_34_4# 2.60fF
C1469 vdd DFFPOSX1_77/a_2_6# 5.17fF
C1470 vdd XOR2X1_50/Y 10.41fF
C1471 vdd XOR2X1_80/a_13_43# 2.11fF
C1472 vdd OAI21X1_0/A 13.20fF
C1473 vdd XNOR2X1_8/a_2_6# 2.29fF
C1474 vdd DFFPOSX1_95/a_2_6# 5.17fF
C1475 XOR2X1_81/A XOR2X1_17/B 2.31fF
C1476 vdd XOR2X1_57/Y 8.55fF
C1477 vdd DFFPOSX1_84/a_2_6# 5.17fF
C1478 vdd INVX2_122/Y 8.35fF
C1479 vdd AOI22X1_94/C 2.68fF
C1480 vdd XNOR2X1_9/A 5.89fF
C1481 vdd BUFX2_7/Y 5.59fF
C1482 XOR2X1_73/a_13_43# vdd 2.11fF
C1483 XOR2X1_29/a_13_43# INVX2_28/Y 2.83fF
C1484 vdd INVX2_110/Y 6.08fF
C1485 vdd AND2X2_9/Y 4.57fF
C1486 vdd XNOR2X1_41/Y 9.19fF
C1487 vdd DFFPOSX1_48/a_22_6# 2.55fF
C1488 DFFPOSX1_55/a_2_6# vdd 5.17fF
C1489 vdd XOR2X1_82/a_2_6# 2.07fF
C1490 XOR2X1_91/A AND2X2_41/a_2_6# 2.51fF
C1491 vdd XOR2X1_61/A 5.38fF
C1492 vdd DFFPOSX1_13/a_22_6# 2.55fF
C1493 XOR2X1_81/a_2_6# XOR2X1_81/A 2.63fF
C1494 vdd NOR2X1_27/Y 4.24fF
C1495 vdd BUFX2_4/Y 34.14fF
C1496 vdd XOR2X1_2/Y 15.82fF
C1497 INVX2_126/Y INVX2_43/Y 2.44fF
C1498 DFFPOSX1_12/a_22_6# vdd 2.55fF
C1499 INVX2_50/Y INVX2_39/A 2.09fF
C1500 vdd HAX1_9/a_2_74# 3.67fF
C1501 vdd INVX2_79/A 2.17fF
C1502 vdd NOR2X1_16/A 11.53fF
C1503 OAI22X1_13/Y vdd 5.30fF
C1504 vdd HAX1_12/YS 5.93fF
C1505 in_inp gnd 2.37fF
C1506 out_MuxData[8] out_MuxData[10] 2.27fF
C1507 vdd HAX1_0/B 5.98fF
C1508 INVX2_87/Y gnd 12.61fF
C1509 vdd XOR2X1_86/a_13_43# 2.11fF
C1510 DFFPOSX1_41/a_2_6# vdd 5.17fF
C1511 AND2X2_26/Y BUFX2_9/Y 2.14fF
C1512 vdd XNOR2X1_6/a_2_6# 2.29fF
C1513 AND2X2_25/Y vdd 3.56fF
C1514 DFFPOSX1_18/a_34_4# vdd 2.60fF
C1515 vdd XOR2X1_60/Y 2.90fF
C1516 vdd XNOR2X1_27/a_2_6# 2.29fF
C1517 vdd DFFPOSX1_9/a_22_6# 2.55fF
C1518 XOR2X1_13/Y gnd 2.32fF
C1519 BUFX2_9/Y INVX2_126/A 2.78fF
C1520 vdd DFFPOSX1_74/a_22_6# 2.55fF
C1521 out_MuxData[8] gnd 12.88fF
C1522 out_MemBData[9] gnd 3.97fF
C1523 vdd XNOR2X1_35/a_2_6# 2.29fF
C1524 vdd OAI21X1_39/C 4.33fF
C1525 vdd DFFPOSX1_5/a_22_6# 2.55fF
C1526 XOR2X1_69/B XOR2X1_38/a_13_43# 3.22fF
C1527 INVX2_104/Y gnd 5.02fF
C1528 INVX2_84/Y gnd 2.68fF
C1529 AOI22X1_74/a_2_54# vdd 2.85fF
C1530 INVX2_82/A vdd 3.15fF
C1531 vdd DFFPOSX1_76/a_22_6# 2.55fF
C1532 XNOR2X1_19/a_2_6# vdd 2.29fF
C1533 AND2X2_39/Y gnd 3.97fF
C1534 vdd NAND2X1_4/Y 4.30fF
C1535 vdd DFFPOSX1_24/a_34_4# 2.60fF
C1536 vdd DFFPOSX1_13/a_34_4# 2.60fF
C1537 con_countWriteout[3] gnd 2.31fF
C1538 XOR2X1_52/a_13_43# INVX2_86/Y 2.57fF
C1539 vdd XNOR2X1_5/a_2_6# 2.29fF
C1540 vdd XOR2X1_82/a_13_43# 2.11fF
C1541 vdd INVX2_40/A 14.81fF
C1542 NOR2X1_0/B out_MuxData[4] 2.27fF
C1543 AOI22X1_48/B OAI21X1_58/Y 2.08fF
C1544 XOR2X1_12/a_2_6# con_countWriteout[8] 2.10fF
C1545 DFFPOSX1_15/a_2_6# vdd 5.17fF
C1546 AND2X2_9/A XOR2X1_21/a_2_6# 2.57fF
C1547 out_MuxData[11] OAI21X1_87/A 3.07fF
C1548 out_state[2] BUFX2_9/Y 2.89fF
C1549 DFFPOSX1_69/a_34_4# vdd 2.60fF
C1550 vdd INVX2_119/Y 5.37fF
C1551 vdd NOR2X1_27/A 4.20fF
C1552 XOR2X1_59/a_2_6# vdd 2.07fF
C1553 vdd XNOR2X1_56/a_2_6# 2.29fF
C1554 vdd NOR2X1_36/Y 3.14fF
C1555 vdd DFFPOSX1_99/a_34_4# 2.60fF
C1556 vdd AOI22X1_89/a_2_54# 2.85fF
C1557 vdd AOI22X1_31/a_2_54# 2.85fF
C1558 vdd BUFX2_7/a_2_6# 2.41fF
C1559 DFFPOSX1_62/a_34_4# INVX2_84/Y 2.45fF
C1560 NOR2X1_3/B vdd 3.85fF
C1561 XOR2X1_69/A XNOR2X1_55/a_2_6# 2.10fF
C1562 vdd AOI22X1_92/a_2_54# 2.85fF
C1563 OAI21X1_45/Y vdd 3.53fF
C1564 vdd OAI21X1_9/Y 2.68fF
C1565 AND2X2_39/B AOI22X1_91/a_2_54# 2.03fF
C1566 XOR2X1_65/A AOI22X1_58/Y 2.53fF
C1567 vdd DFFPOSX1_29/a_22_6# 2.55fF
C1568 vdd DFFPOSX1_82/a_22_6# 2.55fF
C1569 vdd DFFPOSX1_44/a_2_6# 5.17fF
C1570 vdd OAI21X1_31/C 6.25fF
C1571 INVX2_41/Y INVX2_11/Y 2.56fF
C1572 vdd DFFPOSX1_59/a_22_6# 2.55fF
C1573 vdd HAX1_11/YS 3.58fF
C1574 vdd XOR2X1_46/a_2_6# 2.07fF
C1575 vdd XNOR2X1_0/a_2_6# 2.29fF
C1576 vdd XOR2X1_44/Y 4.60fF
C1577 vdd INVX2_118/A 5.53fF
C1578 vdd NOR2X1_16/B 24.74fF
C1579 vdd BUFX2_6/a_2_6# 2.41fF
C1580 vdd AOI22X1_98/a_2_54# 2.85fF
C1581 AND2X2_6/B HAX1_3/YS 2.29fF
C1582 DFFPOSX1_2/a_2_6# vdd 5.17fF
C1583 NOR2X1_8/B XNOR2X1_10/a_2_6# 2.79fF
C1584 DFFPOSX1_57/a_22_6# BUFX2_9/Y 2.71fF
C1585 NOR2X1_40/Y vdd 6.95fF
C1586 DFFPOSX1_62/a_2_6# vdd 5.17fF
C1587 vdd XOR2X1_81/Y 2.92fF
C1588 XOR2X1_55/A AND2X2_23/a_2_6# 2.72fF
C1589 vdd XNOR2X1_54/a_2_6# 2.29fF
C1590 vdd DFFPOSX1_27/a_2_6# 5.04fF
C1591 NOR2X1_23/Y INVX2_92/Y 5.46fF
C1592 vdd DFFPOSX1_94/a_2_6# 5.17fF
C1593 vdd NOR2X1_2/A 3.32fF
C1594 vdd INVX2_76/Y 4.04fF
C1595 XOR2X1_50/B XOR2X1_50/a_13_43# 2.35fF
C1596 vdd DFFPOSX1_42/a_34_4# 2.60fF
C1597 vdd OAI21X1_90/C 8.16fF
C1598 vdd DFFPOSX1_4/a_22_6# 2.55fF
C1599 DFFPOSX1_63/a_22_6# vdd 2.55fF
C1600 vdd INVX2_102/Y 2.35fF
C1601 vdd OR2X1_1/B 5.65fF
C1602 con_loadData gnd 2.22fF
C1603 NOR2X1_12/A XNOR2X1_23/a_12_41# 2.64fF
C1604 XOR2X1_15/a_2_6# vdd 2.07fF
C1605 DFFPOSX1_38/a_22_6# vdd 2.55fF
C1606 INVX2_41/Y DFFPOSX1_13/a_22_6# 2.53fF
C1607 vdd DFFPOSX1_89/a_34_4# 2.60fF
C1608 vdd XOR2X1_24/a_13_43# 2.11fF
C1609 vdd XOR2X1_45/Y 2.09fF
C1610 BUFX2_9/Y INVX2_43/Y 5.47fF
C1611 vdd out_MemBData[7] 9.74fF
C1612 INVX2_86/Y out_MuxData[3] 2.01fF
C1613 AND2X2_18/a_2_6# AND2X2_18/B 2.24fF
C1614 con_countWriteout[6] gnd 3.13fF
C1615 vdd XNOR2X1_28/a_2_6# 2.29fF
C1616 NAND3X1_12/Y DFFPOSX1_25/a_2_6# 2.27fF
C1617 vdd DFFPOSX1_28/a_22_6# 2.55fF
C1618 XOR2X1_50/A out_MuxData[4] 2.67fF
C1619 vdd XNOR2X1_5/Y 3.35fF
C1620 INVX2_57/Y gnd 2.02fF
C1621 BUFX2_10/Y INVX2_84/Y 2.53fF
C1622 INVX2_12/A INVX2_11/A 2.94fF
C1623 XOR2X1_58/Y vdd 4.71fF
C1624 out_MuxData[8] XOR2X1_64/a_2_6# 2.00fF
C1625 XOR2X1_74/a_2_6# out_MuxData[10] 2.01fF
C1626 vdd NOR2X1_47/B 2.41fF
C1627 vdd XOR2X1_1/a_13_43# 2.11fF
C1628 vdd INVX2_69/A 4.93fF
C1629 vdd XOR2X1_56/a_13_43# 2.11fF
C1630 vdd XOR2X1_22/a_13_43# 2.11fF
C1631 vdd AOI22X1_1/a_2_54# 2.85fF
C1632 XOR2X1_69/B XNOR2X1_17/a_2_6# 2.10fF
C1633 XOR2X1_72/a_2_6# vdd 2.07fF
C1634 INVX2_98/Y vdd 8.02fF
C1635 INVX2_82/Y vdd 3.01fF
C1636 BUFX2_10/Y DFFPOSX1_98/a_22_6# 2.31fF
C1637 vdd out_MemBData[8] 14.23fF
C1638 vdd XOR2X1_49/a_13_43# 2.11fF
C1639 vdd AOI22X1_85/a_2_54# 2.85fF
C1640 con_countWriteout[4] vdd 16.58fF
C1641 INVX2_82/A INVX2_99/A 3.19fF
C1642 INVX2_99/Y gnd 2.23fF
C1643 vdd XOR2X1_32/a_2_6# 2.07fF
C1644 vdd XOR2X1_79/Y 3.65fF
C1645 vdd BUFX2_8/Y 11.95fF
C1646 vdd XNOR2X1_14/a_2_6# 2.29fF
C1647 OAI21X1_89/A out_MuxData[8] 2.09fF
C1648 vdd XOR2X1_76/a_2_6# 2.07fF
C1649 INVX2_41/Y vdd 67.97fF
C1650 XNOR2X1_52/a_2_6# XOR2X1_17/B 2.89fF
C1651 XNOR2X1_45/a_2_6# vdd 2.29fF
C1652 vdd AOI22X1_88/C 2.68fF
C1653 vdd INVX2_121/A 2.44fF
C1654 DFFPOSX1_41/a_22_6# vdd 2.55fF
C1655 vdd out_state[0] 9.49fF
C1656 out_MemBData[3] DFFPOSX1_6/a_2_6# 2.15fF
C1657 vdd OAI21X1_78/A 3.91fF
C1658 vdd XOR2X1_78/B 3.03fF
C1659 vdd DFFPOSX1_100/a_2_6# 5.17fF
C1660 vdd DFFPOSX1_30/a_34_4# 2.60fF
C1661 vdd DFFPOSX1_21/a_34_4# 2.60fF
C1662 vdd DFFPOSX1_46/a_34_4# 2.60fF
C1663 vdd INVX2_99/A 8.74fF
C1664 vdd DFFPOSX1_93/a_22_6# 2.55fF
C1665 vdd DFFPOSX1_14/a_22_6# 2.55fF
C1666 INVX2_61/Y BUFX2_4/Y 2.25fF
C1667 BUFX2_8/A vdd 10.17fF
C1668 vdd AND2X2_10/Y 5.82fF
C1669 vdd INVX2_110/A 2.44fF
C1670 AND2X2_9/A vdd 5.00fF
C1671 DFFPOSX1_67/a_22_6# vdd 2.55fF
C1672 AOI22X1_69/B vdd 4.59fF
C1673 vdd AOI22X1_40/a_2_54# 2.85fF
C1674 vdd XOR2X1_24/a_2_6# 2.07fF
C1675 vdd XOR2X1_31/a_2_6# 2.07fF
C1676 vdd XNOR2X1_51/a_2_6# 2.29fF
C1677 vdd XOR2X1_35/a_13_43# 2.11fF
C1678 vdd INVX2_75/A 7.01fF
C1679 vdd NAND3X1_7/A 2.85fF
C1680 vdd AOI21X1_5/Y 3.17fF
C1681 vdd DFFPOSX1_6/a_22_6# 2.55fF
C1682 vdd AOI22X1_29/a_2_54# 2.85fF
C1683 XOR2X1_74/Y vdd 4.89fF
C1684 XOR2X1_10/a_2_6# vdd 2.07fF
C1685 XNOR2X1_29/a_2_6# INVX2_86/Y 2.10fF
C1686 vdd INVX2_133/Y 4.83fF
C1687 out_temp_addNum[1] gnd 6.67fF
C1688 vdd XOR2X1_0/a_2_6# 2.07fF
C1689 vdd XNOR2X1_7/A 5.05fF
C1690 vdd HAX1_6/B 5.32fF
C1691 XOR2X1_37/B XOR2X1_37/a_13_43# 2.64fF
C1692 out_MuxData[8] XOR2X1_64/Y 2.25fF
C1693 XNOR2X1_16/a_2_6# vdd 2.29fF
C1694 DFFPOSX1_6/a_34_4# vdd 2.60fF
C1695 out_MuxData[7] out_MuxData[8] 2.87fF
C1696 vdd XOR2X1_47/a_2_6# 2.07fF
C1697 vdd XOR2X1_21/Y 5.38fF
C1698 vdd DFFPOSX1_9/a_2_6# 5.17fF
C1699 vdd XNOR2X1_7/a_2_6# 2.29fF
C1700 vdd OAI21X1_50/B 5.19fF
C1701 vdd DFFPOSX1_16/a_2_6# 5.17fF
C1702 XNOR2X1_3/a_2_6# OAI21X1_5/Y 2.10fF
C1703 vdd XOR2X1_6/a_13_43# 2.11fF
C1704 vdd XOR2X1_89/a_2_6# 2.07fF
C1705 BUFX2_10/Y DFFPOSX1_86/a_22_6# 2.25fF
C1706 XNOR2X1_31/a_2_6# XOR2X1_81/A 3.98fF
C1707 AND2X2_25/a_2_6# INVX2_72/Y 2.10fF
C1708 BUFX2_10/a_2_6# vdd 2.41fF
C1709 con_count[6] BUFX2_9/Y 3.61fF
C1710 XNOR2X1_21/a_12_41# XOR2X1_43/Y 2.91fF
C1711 vdd NOR2X1_14/Y 5.83fF
C1712 DFFPOSX1_41/a_34_4# out_MuxData[10] 2.22fF
C1713 vdd INVX2_61/Y 55.99fF
C1714 vdd XOR2X1_60/a_2_6# 2.07fF
C1715 vdd DFFPOSX1_77/a_22_6# 2.55fF
C1716 OAI22X1_9/Y BUFX2_11/Y 2.55fF
C1717 vdd INVX2_44/A 8.07fF
C1718 vdd INVX2_85/Y 8.30fF
C1719 vdd XOR2X1_87/a_13_43# 2.11fF
C1720 BUFX2_10/Y DFFPOSX1_58/a_22_6# 2.31fF
C1721 AOI22X1_48/a_2_54# INVX2_92/Y 2.18fF
C1722 out_MuxData[11] vdd 54.60fF
C1723 vdd NAND3X1_25/B 7.80fF
C1724 out_MuxData[9] XOR2X1_17/B 2.10fF
C1725 vdd NOR2X1_22/Y 20.53fF
C1726 out_MuxData[1] out_MuxData[2] 2.31fF
C1727 HAX1_7/YS vdd 3.19fF
C1728 DFFPOSX1_69/a_2_6# vdd 5.17fF
C1729 AOI22X1_27/a_2_54# vdd 2.85fF
C1730 vdd AOI22X1_51/B 6.96fF
C1731 DFFPOSX1_23/a_34_4# vdd 2.60fF
C1732 AND2X2_20/A vdd 10.66fF
C1733 vdd XOR2X1_64/a_13_43# 2.11fF
C1734 con_count[5] gnd 3.46fF
C1735 vdd AND2X2_21/Y 11.74fF
C1736 vdd AOI22X1_0/C 2.68fF
C1737 vdd DFFPOSX1_99/a_2_6# 5.17fF
C1738 vdd XOR2X1_90/a_2_6# 2.07fF
C1739 INVX2_46/A con_restart 2.25fF
C1740 INVX2_46/A INVX2_59/Y 2.93fF
C1741 NOR2X1_14/B XNOR2X1_24/a_2_6# 2.10fF
C1742 vdd OR2X1_1/Y 3.63fF
C1743 AND2X2_6/B BUFX2_5/Y 2.06fF
C1744 vdd DFFPOSX1_90/a_22_6# 2.55fF
C1745 NOR2X1_46/B NOR2X1_46/Y 2.13fF
C1746 gnd AND2X2_4/A 5.91fF
C1747 AOI21X1_4/Y vdd 2.76fF
C1748 vdd NAND3X1_22/B 8.38fF
C1749 vdd INVX2_64/Y 4.15fF
C1750 out_MuxData[1] XOR2X1_79/a_2_6# 2.37fF
C1751 vdd XOR2X1_5/a_2_6# 2.07fF
C1752 vdd XOR2X1_48/Y 4.19fF
C1753 INVX2_43/Y INVX2_126/A 3.02fF
C1754 INVX2_28/Y gnd 7.62fF
C1755 vdd INVX2_27/Y 3.72fF
C1756 vdd XOR2X1_85/a_13_43# 2.11fF
C1757 vdd DFFPOSX1_54/a_34_4# 2.60fF
C1758 vdd XNOR2X1_55/a_2_6# 2.29fF
C1759 INVX2_59/Y out_MuxData[15] 3.52fF
C1760 vdd AOI22X1_2/a_2_54# 2.85fF
C1761 NAND2X1_8/Y vdd 8.34fF
C1762 OAI21X1_65/C vdd 4.00fF
C1763 INVX2_11/Y INVX2_11/A 2.48fF
C1764 BUFX2_10/Y DFFPOSX1_83/a_22_6# 2.25fF
C1765 vdd DFFPOSX1_59/a_2_6# 5.17fF
C1766 vdd NAND3X1_8/Y 7.72fF
C1767 vdd AND2X2_14/A 10.51fF
C1768 vdd XNOR2X1_27/A 5.74fF
C1769 vdd INVX2_51/A 19.86fF
C1770 vdd XOR2X1_89/B 5.84fF
C1771 BUFX2_11/Y OR2X2_0/Y 2.47fF
C1772 INVX2_16/Y XNOR2X1_13/a_2_6# 2.64fF
C1773 INVX2_116/A INVX2_126/A 2.00fF
C1774 vdd DFFPOSX1_18/a_22_6# 2.55fF
C1775 vdd XOR2X1_58/A 5.72fF
C1776 vdd NAND3X1_2/Y 9.34fF
C1777 vdd INVX2_127/Y 3.11fF
C1778 vdd AOI22X1_11/a_2_54# 2.85fF
C1779 vdd XOR2X1_21/a_13_43# 2.11fF
C1780 gnd AND2X2_18/A 2.03fF
C1781 AND2X2_6/B gnd 4.11fF
C1782 AND2X2_21/B vdd 5.14fF
C1783 vdd XOR2X1_9/Y 2.59fF
C1784 vdd XOR2X1_75/a_2_6# 2.07fF
C1785 vdd DFFPOSX1_78/a_22_6# 2.55fF
C1786 vdd DFFPOSX1_89/a_2_6# 5.17fF
C1787 DFFPOSX1_35/a_2_6# vdd 5.17fF
C1788 DFFPOSX1_40/a_2_6# vdd 5.17fF
C1789 XOR2X1_77/a_13_43# XOR2X1_17/B 3.65fF
C1790 vdd XOR2X1_28/B 3.79fF
C1791 vdd con_countWriteout[2] 19.36fF
C1792 INVX2_41/Y DFFPOSX1_6/a_22_6# 2.09fF
C1793 vdd NAND3X1_34/B 9.32fF
C1794 vdd OAI21X1_32/C 7.71fF
C1795 INVX2_59/A out_MemBData[15] 2.55fF
C1796 vdd XOR2X1_26/a_13_43# 2.11fF
C1797 vdd AOI22X1_94/a_2_54# 2.85fF
C1798 vdd DFFPOSX1_96/a_22_6# 2.55fF
C1799 vdd DFFPOSX1_53/a_34_4# 2.60fF
C1800 vdd XOR2X1_18/a_2_6# 2.07fF
C1801 con_countWriteout[7] BUFX2_5/Y 2.23fF
C1802 INVX2_38/Y vdd 5.49fF
C1803 AOI22X1_24/a_2_54# vdd 2.85fF
C1804 vdd HAX1_10/a_2_74# 3.67fF
C1805 vdd NOR2X1_44/A 2.22fF
C1806 vdd DFFPOSX1_80/a_2_6# 5.17fF
C1807 XOR2X1_62/a_13_43# vdd 2.11fF
C1808 out_MemBData[13] NOR2X1_23/Y 2.46fF
C1809 vdd DFFPOSX1_27/a_22_6# 2.55fF
C1810 INVX2_16/Y AND2X2_9/B 2.04fF
C1811 vdd XNOR2X1_26/a_2_6# 2.29fF
C1812 INVX2_80/A INVX2_126/A 3.12fF
C1813 OAI21X1_35/B gnd 2.00fF
C1814 vdd XOR2X1_63/Y 3.40fF
C1815 vdd XOR2X1_82/Y 3.33fF
C1816 vdd out_MuxData[14] 35.56fF
C1817 vdd AOI22X1_48/B 10.53fF
C1818 NAND3X1_27/B OAI21X1_68/B 2.49fF
C1819 out_MuxData[8] out_MuxData[9] 2.70fF
C1820 vdd OAI21X1_79/C 7.92fF
C1821 vdd XOR2X1_3/a_2_6# 2.07fF
C1822 vdd NAND3X1_0/Y 6.91fF
C1823 vdd INVX2_86/Y 21.99fF
C1824 vdd OAI22X1_5/Y 3.02fF
C1825 vdd OAI21X1_89/C 9.28fF
C1826 out_MemBData[5] OR2X2_0/Y 2.71fF
C1827 INVX2_35/Y vdd 4.11fF
C1828 AND2X2_28/B OAI22X1_6/C 2.03fF
C1829 INVX2_56/Y BUFX2_2/Y 2.60fF
C1830 con_count[7] vdd 7.35fF
C1831 XOR2X1_27/A vdd 3.66fF
C1832 XOR2X1_51/Y AND2X2_17/Y 2.91fF
C1833 INVX2_52/Y gnd 2.63fF
C1834 XNOR2X1_41/a_2_6# vdd 2.29fF
C1835 vdd INVX2_40/Y 8.54fF
C1836 INVX2_43/Y INVX2_53/A 2.29fF
C1837 vdd AOI22X1_2/C 3.77fF
C1838 vdd in_reset 6.55fF
C1839 vdd XOR2X1_37/B 4.23fF
C1840 INVX2_126/Y gnd 9.91fF
C1841 vdd INVX2_36/Y 3.04fF
C1842 AND2X2_9/B out_MuxData[6] 2.18fF
C1843 INVX2_89/A INVX2_126/A 2.22fF
C1844 BUFX2_10/Y DFFPOSX1_70/a_22_6# 2.31fF
C1845 vdd XOR2X1_76/a_13_43# 2.11fF
C1846 NOR2X1_32/Y vdd 6.08fF
C1847 vdd DFFPOSX1_81/a_22_6# 2.55fF
C1848 vdd DFFPOSX1_88/a_22_6# 2.55fF
C1849 DFFPOSX1_66/a_22_6# vdd 2.55fF
C1850 con_countWriteout[8] vdd 10.47fF
C1851 vdd DFFPOSX1_45/a_22_6# 2.55fF
C1852 vdd XNOR2X1_9/a_2_6# 2.29fF
C1853 vdd AND2X2_8/Y 2.82fF
C1854 vdd AOI21X1_7/A 2.86fF
C1855 INVX2_41/Y OR2X1_1/Y 2.25fF
C1856 vdd INVX2_11/A 43.43fF
C1857 vdd XOR2X1_78/a_2_6# 2.07fF
C1858 vdd AOI22X1_20/a_2_54# 2.85fF
C1859 vdd XOR2X1_36/a_13_43# 2.11fF
C1860 vdd DFFPOSX1_93/a_34_4# 2.60fF
C1861 XOR2X1_69/B out_MuxData[10] 2.38fF
C1862 OAI21X1_89/A XOR2X1_91/A 2.23fF
C1863 XOR2X1_53/Y vdd 3.00fF
C1864 vdd HAX1_10/B 3.34fF
C1865 vdd AND2X2_20/B 2.52fF
C1866 vdd DFFPOSX1_86/a_34_4# 2.60fF
C1867 vdd AOI22X1_58/Y 9.60fF
C1868 XOR2X1_33/a_2_6# XOR2X1_33/A 2.57fF
C1869 DFFPOSX1_67/a_34_4# vdd 2.60fF
C1870 vdd DFFPOSX1_48/a_34_4# 2.60fF
C1871 XOR2X1_59/Y vdd 2.57fF
C1872 INVX2_88/Y vdd 5.90fF
C1873 BUFX2_9/Y INVX2_72/Y 3.09fF
C1874 vdd XOR2X1_4/a_2_6# 2.07fF
C1875 vdd INVX2_25/A 19.54fF
C1876 in_clka gnd 3.49fF
C1877 vdd XNOR2X1_20/a_2_6# 2.29fF
C1878 XOR2X1_69/B gnd 3.51fF
C1879 vdd DFFPOSX1_75/a_22_6# 2.55fF
C1880 vdd XOR2X1_45/a_13_43# 2.11fF
C1881 vdd INVX2_75/Y 30.48fF
C1882 con_countWriteout[1] Gnd 23.36fF
C1883 con_countWriteout[3] Gnd 8.55fF
C1884 con_countWriteout[4] Gnd 26.48fF
C1885 gnd Gnd 5668.64fF
C1886 con_countWriteout[7] Gnd 25.75fF
C1887 BUFX2_5/Y Gnd 94.55fF
C1888 out_MemBData[3] Gnd 19.86fF
C1889 NAND3X1_2/Y Gnd 5.55fF
C1890 INVX2_6/A Gnd 8.87fF
C1891 vdd Gnd 23516.19fF
C1892 out_MuxData[12] Gnd 92.16fF
C1893 DFFPOSX1_0/a_66_6# Gnd 2.23fF
C1894 DFFPOSX1_0/a_2_6# Gnd 3.02fF
C1895 INVX2_1/Y Gnd 8.63fF
C1896 DFFPOSX1_1/a_66_6# Gnd 2.23fF
C1897 AOI22X1_0/C Gnd 8.97fF
C1898 DFFPOSX1_1/a_2_6# Gnd 3.02fF
C1899 AND2X2_0/Y Gnd 8.85fF
C1900 AND2X2_0/a_2_6# Gnd 2.37fF
C1901 DFFPOSX1_2/a_66_6# Gnd 2.23fF
C1902 AOI22X1_1/C Gnd 11.99fF
C1903 DFFPOSX1_2/a_2_6# Gnd 3.02fF
C1904 AND2X2_1/Y Gnd 2.85fF
C1905 AND2X2_1/a_2_6# Gnd 2.37fF
C1906 AND2X2_2/a_2_6# Gnd 2.37fF
C1907 DFFPOSX1_3/a_66_6# Gnd 2.23fF
C1908 con_countWriteout[5] Gnd 21.95fF
C1909 DFFPOSX1_3/a_2_6# Gnd 3.02fF
C1910 INVX2_0/Y Gnd 8.79fF
C1911 AND2X2_3/a_2_6# Gnd 2.37fF
C1912 DFFPOSX1_5/a_66_6# Gnd 2.23fF
C1913 AOI22X1_3/C Gnd 8.53fF
C1914 DFFPOSX1_5/a_2_6# Gnd 3.02fF
C1915 AND2X2_3/Y Gnd 9.22fF
C1916 DFFPOSX1_6/a_66_6# Gnd 2.23fF
C1917 DFFPOSX1_6/a_2_6# Gnd 3.02fF
C1918 INVX2_2/Y Gnd 5.82fF
C1919 XOR2X1_0/a_2_6# Gnd 3.50fF
C1920 XOR2X1_0/a_13_43# Gnd 3.05fF
C1921 XOR2X1_0/A Gnd 3.12fF
C1922 INVX2_3/Y Gnd 9.72fF
C1923 XNOR2X1_0/a_2_6# Gnd 2.31fF
C1924 XNOR2X1_0/a_12_41# Gnd 3.38fF
C1925 AND2X2_4/a_2_6# Gnd 2.37fF
C1926 XNOR2X1_0/A Gnd 10.06fF
C1927 XOR2X1_1/B Gnd 12.96fF
C1928 OAI21X1_2/C Gnd 10.19fF
C1929 AND2X2_4/A Gnd 25.07fF
C1930 NAND3X1_0/Y Gnd 7.63fF
C1931 OAI21X1_2/A Gnd 3.56fF
C1932 XOR2X1_2/a_2_6# Gnd 3.50fF
C1933 XOR2X1_2/a_13_43# Gnd 3.05fF
C1934 XOR2X1_2/A Gnd 3.06fF
C1935 XOR2X1_3/Y Gnd 17.11fF
C1936 XOR2X1_3/a_2_6# Gnd 3.50fF
C1937 XOR2X1_3/a_13_43# Gnd 3.05fF
C1938 XOR2X1_2/B Gnd 6.33fF
C1939 INVX2_4/Y Gnd 3.66fF
C1940 INVX2_4/A Gnd 5.49fF
C1941 AND2X2_5/A Gnd 14.50fF
C1942 XNOR2X1_2/a_2_6# Gnd 2.31fF
C1943 XNOR2X1_2/a_12_41# Gnd 3.38fF
C1944 NOR2X1_2/B Gnd 14.58fF
C1945 NOR2X1_2/A Gnd 12.10fF
C1946 NOR2X1_2/Y Gnd 10.50fF
C1947 XOR2X1_7/a_2_6# Gnd 3.50fF
C1948 XOR2X1_7/a_13_43# Gnd 3.05fF
C1949 XOR2X1_7/A Gnd 5.11fF
C1950 NAND3X1_1/Y Gnd 4.82fF
C1951 NAND3X1_1/B Gnd 12.47fF
C1952 INVX2_6/Y Gnd 15.79fF
C1953 OAI21X1_4/A Gnd 15.44fF
C1954 XOR2X1_8/a_2_6# Gnd 3.50fF
C1955 XOR2X1_8/a_13_43# Gnd 3.05fF
C1956 NAND2X1_3/A Gnd 10.33fF
C1957 XOR2X1_8/Y Gnd 9.18fF
C1958 out_MuxData[6] Gnd 3.86fF
C1959 out_MuxData[2] Gnd 47.99fF
C1960 NAND3X1_4/B Gnd 7.54fF
C1961 OAI21X1_6/B Gnd 20.30fF
C1962 out_MemBData[1] Gnd 21.47fF
C1963 INVX2_11/A Gnd 13.76fF
C1964 INVX2_28/Y Gnd 17.58fF
C1965 INVX2_1/A Gnd 8.04fF
C1966 HAX1_0/YS Gnd 3.74fF
C1967 HAX1_0/YC Gnd 3.52fF
C1968 HAX1_0/a_41_74# Gnd 2.55fF
C1969 HAX1_0/a_2_74# Gnd 2.94fF
C1970 OR2X1_1/B Gnd 6.26fF
C1971 OR2X1_0/a_2_54# Gnd 2.68fF
C1972 con_countWriteout[8] Gnd 22.53fF
C1973 INVX2_9/A Gnd 7.77fF
C1974 HAX1_1/YS Gnd 9.02fF
C1975 HAX1_0/B Gnd 6.41fF
C1976 HAX1_1/a_41_74# Gnd 2.55fF
C1977 HAX1_1/a_2_74# Gnd 2.94fF
C1978 con_countWriteout[6] Gnd 18.84fF
C1979 HAX1_1/B Gnd 6.24fF
C1980 HAX1_2/a_41_74# Gnd 2.55fF
C1981 HAX1_2/a_2_74# Gnd 2.94fF
C1982 DFFPOSX1_4/a_66_6# Gnd 2.23fF
C1983 DFFPOSX1_4/a_2_6# Gnd 3.02fF
C1984 INVX2_0/A Gnd 4.08fF
C1985 AOI22X1_2/C Gnd 9.23fF
C1986 HAX1_3/YS Gnd 8.60fF
C1987 HAX1_2/B Gnd 6.29fF
C1988 HAX1_3/a_41_74# Gnd 2.55fF
C1989 HAX1_3/a_2_74# Gnd 2.94fF
C1990 HAX1_3/B Gnd 10.02fF
C1991 INVX2_11/Y Gnd 6.42fF
C1992 INVX2_2/A Gnd 7.67fF
C1993 DFFPOSX1_7/a_66_6# Gnd 2.23fF
C1994 DFFPOSX1_7/a_2_6# Gnd 3.02fF
C1995 INVX2_15/Y Gnd 8.28fF
C1996 INVX2_41/Y Gnd 86.58fF
C1997 XNOR2X1_7/A Gnd 11.16fF
C1998 NAND3X1_2/B Gnd 8.16fF
C1999 OAI21X1_0/A Gnd 3.77fF
C2000 INVX2_3/A Gnd 8.13fF
C2001 XOR2X1_0/B Gnd 16.98fF
C2002 NOR2X1_0/B Gnd 11.44fF
C2003 XOR2X1_1/a_2_6# Gnd 3.50fF
C2004 XOR2X1_1/a_13_43# Gnd 3.05fF
C2005 XNOR2X1_1/a_2_6# Gnd 2.31fF
C2006 XNOR2X1_1/a_12_41# Gnd 3.38fF
C2007 NOR2X1_0/A Gnd 13.75fF
C2008 XOR2X1_15/B Gnd 7.77fF
C2009 out_MuxData[14] Gnd 52.85fF
C2010 XOR2X1_4/Y Gnd 10.09fF
C2011 out_MuxData[10] Gnd 47.43fF
C2012 XOR2X1_4/a_2_6# Gnd 3.50fF
C2013 XOR2X1_4/a_13_43# Gnd 3.05fF
C2014 out_MuxData[4] Gnd 49.54fF
C2015 XOR2X1_5/a_2_6# Gnd 3.50fF
C2016 XOR2X1_5/a_13_43# Gnd 3.05fF
C2017 out_MuxData[5] Gnd 22.54fF
C2018 XOR2X1_5/A Gnd 10.73fF
C2019 XOR2X1_6/a_2_6# Gnd 3.50fF
C2020 XOR2X1_6/a_13_43# Gnd 3.05fF
C2021 XOR2X1_6/A Gnd 8.79fF
C2022 INVX2_5/A Gnd 30.11fF
C2023 out_MuxData[15] Gnd 50.12fF
C2024 XOR2X1_9/Y Gnd 13.84fF
C2025 XOR2X1_9/a_2_6# Gnd 3.50fF
C2026 XOR2X1_9/a_13_43# Gnd 3.05fF
C2027 XOR2X1_9/B Gnd 9.74fF
C2028 XOR2X1_19/Y Gnd 13.56fF
C2029 XOR2X1_10/a_2_6# Gnd 3.50fF
C2030 XOR2X1_10/a_13_43# Gnd 3.05fF
C2031 XOR2X1_11/a_2_6# Gnd 3.50fF
C2032 XOR2X1_11/a_13_43# Gnd 3.05fF
C2033 AND2X2_5/a_2_6# Gnd 2.37fF
C2034 AND2X2_5/B Gnd 11.61fF
C2035 XNOR2X1_3/Y Gnd 5.00fF
C2036 AND2X2_5/Y Gnd 3.57fF
C2037 XNOR2X1_3/a_2_6# Gnd 2.31fF
C2038 XNOR2X1_3/a_12_41# Gnd 3.38fF
C2039 OAI21X1_5/Y Gnd 8.44fF
C2040 AND2X2_9/B Gnd 14.38fF
C2041 XNOR2X1_4/a_2_6# Gnd 2.31fF
C2042 XNOR2X1_4/a_12_41# Gnd 3.38fF
C2043 INVX2_16/Y Gnd 41.90fF
C2044 XNOR2X1_5/Y Gnd 9.30fF
C2045 XNOR2X1_5/a_2_6# Gnd 2.31fF
C2046 XNOR2X1_5/a_12_41# Gnd 3.38fF
C2047 XNOR2X1_5/A Gnd 7.52fF
C2048 NAND2X1_5/Y Gnd 16.73fF
C2049 INVX2_17/Y Gnd 29.55fF
C2050 XOR2X1_17/B Gnd 36.39fF
C2051 DFFPOSX1_8/a_66_6# Gnd 2.23fF
C2052 DFFPOSX1_8/a_2_6# Gnd 3.02fF
C2053 INVX2_7/Y Gnd 8.11fF
C2054 AOI22X1_9/C Gnd 9.73fF
C2055 AND2X2_6/Y Gnd 8.77fF
C2056 AND2X2_6/a_2_6# Gnd 2.37fF
C2057 AND2X2_6/A Gnd 3.89fF
C2058 XOR2X1_12/a_2_6# Gnd 3.50fF
C2059 XOR2X1_12/a_13_43# Gnd 3.05fF
C2060 DFFPOSX1_10/a_66_6# Gnd 2.23fF
C2061 DFFPOSX1_10/a_2_6# Gnd 3.02fF
C2062 INVX2_9/Y Gnd 8.03fF
C2063 OR2X1_1/a_2_54# Gnd 2.68fF
C2064 OAI21X1_8/Y Gnd 7.48fF
C2065 OR2X1_1/Y Gnd 7.40fF
C2066 OAI21X1_9/Y Gnd 10.04fF
C2067 INVX2_13/Y Gnd 5.18fF
C2068 HAX1_4/YS Gnd 8.22fF
C2069 HAX1_4/a_41_74# Gnd 2.55fF
C2070 HAX1_4/a_2_74# Gnd 2.94fF
C2071 HAX1_4/B Gnd 3.53fF
C2072 INVX2_14/Y Gnd 2.24fF
C2073 AOI22X1_10/C Gnd 8.98fF
C2074 XOR2X1_13/Y Gnd 2.79fF
C2075 XOR2X1_13/a_2_6# Gnd 3.50fF
C2076 XOR2X1_13/a_13_43# Gnd 3.05fF
C2077 AND2X2_8/A Gnd 11.81fF
C2078 XNOR2X1_6/a_2_6# Gnd 2.31fF
C2079 XNOR2X1_6/a_12_41# Gnd 3.38fF
C2080 XOR2X1_14/a_2_6# Gnd 3.50fF
C2081 XOR2X1_14/a_13_43# Gnd 3.05fF
C2082 XNOR2X1_6/B Gnd 10.11fF
C2083 XOR2X1_14/B Gnd 8.77fF
C2084 XOR2X1_15/a_2_6# Gnd 3.50fF
C2085 XOR2X1_15/a_13_43# Gnd 3.05fF
C2086 XOR2X1_16/a_2_6# Gnd 3.50fF
C2087 XOR2X1_16/a_13_43# Gnd 3.05fF
C2088 XOR2X1_18/B Gnd 5.56fF
C2089 XOR2X1_17/a_2_6# Gnd 3.50fF
C2090 XOR2X1_17/a_13_43# Gnd 3.05fF
C2091 out_MuxData[8] Gnd 28.83fF
C2092 XNOR2X1_9/a_2_6# Gnd 2.31fF
C2093 XNOR2X1_9/a_12_41# Gnd 3.38fF
C2094 XNOR2X1_9/A Gnd 26.51fF
C2095 XOR2X1_19/a_2_6# Gnd 3.50fF
C2096 XOR2X1_19/a_13_43# Gnd 3.05fF
C2097 NAND3X1_16/B Gnd 7.18fF
C2098 INVX2_26/Y Gnd 23.43fF
C2099 INVX2_25/Y Gnd 18.75fF
C2100 XOR2X1_30/Y Gnd 13.51fF
C2101 XOR2X1_20/a_2_6# Gnd 3.50fF
C2102 XOR2X1_20/a_13_43# Gnd 3.05fF
C2103 XOR2X1_21/Y Gnd 6.39fF
C2104 XOR2X1_21/a_2_6# Gnd 3.50fF
C2105 XOR2X1_21/a_13_43# Gnd 3.05fF
C2106 AND2X2_9/a_2_6# Gnd 2.37fF
C2107 XOR2X1_22/a_2_6# Gnd 3.50fF
C2108 XOR2X1_22/a_13_43# Gnd 3.05fF
C2109 AND2X2_9/A Gnd 5.52fF
C2110 XOR2X1_24/A Gnd 12.81fF
C2111 AOI21X1_2/Y Gnd 8.72fF
C2112 INVX2_10/A Gnd 2.37fF
C2113 NAND2X1_4/A Gnd 19.01fF
C2114 out_MuxData[13] Gnd 61.94fF
C2115 in_run Gnd 10.88fF
C2116 INVX2_19/A Gnd 16.62fF
C2117 NAND2X1_6/Y Gnd 6.93fF
C2118 INVX2_8/Y Gnd 4.95fF
C2119 DFFPOSX1_9/a_66_6# Gnd 2.23fF
C2120 DFFPOSX1_9/a_2_6# Gnd 3.02fF
C2121 OAI21X1_7/Y Gnd 8.30fF
C2122 AOI21X1_2/B Gnd 2.40fF
C2123 in_wai Gnd 10.63fF
C2124 DFFPOSX1_11/a_66_6# Gnd 2.23fF
C2125 DFFPOSX1_11/a_2_6# Gnd 3.02fF
C2126 INVX2_12/Y Gnd 11.66fF
C2127 INVX2_12/A Gnd 5.52fF
C2128 AND2X2_7/a_2_6# Gnd 2.37fF
C2129 DFFPOSX1_12/a_66_6# Gnd 2.23fF
C2130 DFFPOSX1_12/a_2_6# Gnd 3.02fF
C2131 AND2X2_7/Y Gnd 10.14fF
C2132 DFFPOSX1_13/a_66_6# Gnd 2.23fF
C2133 con_countWriteout[2] Gnd 16.67fF
C2134 DFFPOSX1_13/a_2_6# Gnd 3.02fF
C2135 INVX2_24/Y Gnd 9.36fF
C2136 AND2X2_8/a_2_6# Gnd 2.37fF
C2137 XNOR2X1_7/Y Gnd 4.89fF
C2138 AND2X2_8/Y Gnd 8.94fF
C2139 XNOR2X1_7/a_2_6# Gnd 2.31fF
C2140 XNOR2X1_7/a_12_41# Gnd 3.38fF
C2141 AND2X2_14/Y Gnd 7.15fF
C2142 XNOR2X1_8/a_2_6# Gnd 2.31fF
C2143 XNOR2X1_8/a_12_41# Gnd 3.38fF
C2144 XNOR2X1_8/A Gnd 7.52fF
C2145 NAND2X1_4/Y Gnd 12.23fF
C2146 XOR2X1_27/A Gnd 6.35fF
C2147 NAND3X1_3/Y Gnd 4.12fF
C2148 XOR2X1_18/a_2_6# Gnd 3.50fF
C2149 XOR2X1_18/a_13_43# Gnd 3.05fF
C2150 NAND2X1_4/B Gnd 7.14fF
C2151 NOR2X1_8/A Gnd 15.53fF
C2152 XNOR2X1_10/a_2_6# Gnd 2.31fF
C2153 XNOR2X1_10/a_12_41# Gnd 3.38fF
C2154 NOR2X1_8/B Gnd 12.74fF
C2155 out_MuxData[7] Gnd 41.61fF
C2156 AND2X2_17/A Gnd 10.37fF
C2157 XOR2X1_23/a_2_6# Gnd 3.50fF
C2158 XOR2X1_23/a_13_43# Gnd 3.05fF
C2159 XOR2X1_22/A Gnd 4.91fF
C2160 XOR2X1_23/A Gnd 7.38fF
C2161 XOR2X1_24/a_2_6# Gnd 3.50fF
C2162 XOR2X1_24/a_13_43# Gnd 3.05fF
C2163 NOR2X1_3/Y Gnd 3.70fF
C2164 INVX2_30/Y Gnd 8.09fF
C2165 NOR2X1_3/B Gnd 13.15fF
C2166 XOR2X1_25/a_2_6# Gnd 3.50fF
C2167 XOR2X1_25/a_13_43# Gnd 3.05fF
C2168 INVX2_30/A Gnd 7.05fF
C2169 INVX2_27/Y Gnd 20.10fF
C2170 INVX2_20/Y Gnd 7.58fF
C2171 INVX2_18/Y Gnd 4.84fF
C2172 NAND3X1_6/Y Gnd 7.54fF
C2173 NOR2X1_4/Y Gnd 5.72fF
C2174 INVX2_21/Y Gnd 10.46fF
C2175 con_loseSig Gnd 18.57fF
C2176 INVX2_21/A Gnd 10.89fF
C2177 OAI21X1_28/A Gnd 13.01fF
C2178 INVX2_22/Y Gnd 12.51fF
C2179 AND2X2_10/Y Gnd 8.16fF
C2180 AND2X2_10/a_2_6# Gnd 2.37fF
C2181 AOI22X1_18/C Gnd 8.88fF
C2182 HAX1_5/YS Gnd 8.07fF
C2183 HAX1_5/a_41_74# Gnd 2.55fF
C2184 HAX1_5/a_2_74# Gnd 2.94fF
C2185 con_countWriteout[0] Gnd 35.18fF
C2186 HAX1_6/YS Gnd 5.17fF
C2187 HAX1_6/a_41_74# Gnd 2.55fF
C2188 HAX1_6/a_2_74# Gnd 2.94fF
C2189 HAX1_6/B Gnd 12.05fF
C2190 AND2X2_11/Y Gnd 12.16fF
C2191 AND2X2_11/a_2_6# Gnd 2.37fF
C2192 INVX2_24/A Gnd 4.38fF
C2193 AOI22X1_19/C Gnd 6.72fF
C2194 NAND3X1_7/A Gnd 6.31fF
C2195 NOR2X1_41/B Gnd 13.36fF
C2196 AND2X2_13/a_2_6# Gnd 2.37fF
C2197 AND2X2_13/B Gnd 7.38fF
C2198 AND2X2_14/a_2_6# Gnd 2.37fF
C2199 XOR2X1_26/a_2_6# Gnd 3.50fF
C2200 XOR2X1_26/a_13_43# Gnd 3.05fF
C2201 NAND3X1_3/C Gnd 19.65fF
C2202 XNOR2X1_12/a_2_6# Gnd 2.31fF
C2203 XNOR2X1_12/a_12_41# Gnd 3.38fF
C2204 XOR2X1_35/Y Gnd 10.88fF
C2205 out_MuxData[11] Gnd 46.06fF
C2206 XNOR2X1_13/a_2_6# Gnd 2.31fF
C2207 XNOR2X1_13/a_12_41# Gnd 3.38fF
C2208 XOR2X1_28/Y Gnd 8.93fF
C2209 XOR2X1_28/a_2_6# Gnd 3.50fF
C2210 XOR2X1_28/a_13_43# Gnd 3.05fF
C2211 NAND3X1_8/B Gnd 8.24fF
C2212 XOR2X1_30/a_2_6# Gnd 3.50fF
C2213 XOR2X1_30/a_13_43# Gnd 3.05fF
C2214 out_MuxData[0] Gnd 41.89fF
C2215 XNOR2X1_15/a_2_6# Gnd 2.31fF
C2216 XNOR2X1_15/a_12_41# Gnd 3.38fF
C2217 XNOR2X1_22/A Gnd 13.52fF
C2218 OAI22X1_6/C Gnd 51.87fF
C2219 NAND2X1_8/Y Gnd 10.56fF
C2220 in_inp Gnd 15.20fF
C2221 NOR2X1_5/Y Gnd 2.55fF
C2222 OAI21X1_18/Y Gnd 11.02fF
C2223 con_restart Gnd 75.39fF
C2224 XOR2X1_33/Y Gnd 5.89fF
C2225 AND2X2_15/Y Gnd 3.49fF
C2226 XOR2X1_28/B Gnd 12.79fF
C2227 XNOR2X1_19/A Gnd 4.52fF
C2228 INVX2_19/Y Gnd 6.94fF
C2229 out_state[1] Gnd 25.64fF
C2230 out_state[2] Gnd 35.32fF
C2231 AOI21X1_4/C Gnd 8.11fF
C2232 DFFPOSX1_14/a_66_6# Gnd 2.23fF
C2233 DFFPOSX1_14/a_2_6# Gnd 3.02fF
C2234 AND2X2_12/Y Gnd 10.11fF
C2235 AND2X2_12/a_2_6# Gnd 2.37fF
C2236 DFFPOSX1_15/a_66_6# Gnd 2.23fF
C2237 DFFPOSX1_15/a_2_6# Gnd 3.02fF
C2238 BUFX2_9/Y Gnd 76.04fF
C2239 INVX2_25/A Gnd 18.18fF
C2240 OAI21X1_30/C Gnd 4.73fF
C2241 NOR2X1_6/Y Gnd 4.12fF
C2242 OAI21X1_31/C Gnd 7.89fF
C2243 AND2X2_19/Y Gnd 53.76fF
C2244 NOR2X1_7/Y Gnd 6.80fF
C2245 NAND3X1_7/Y Gnd 17.22fF
C2246 NAND3X1_7/B Gnd 6.84fF
C2247 AND2X2_13/A Gnd 8.47fF
C2248 AOI22X1_23/A Gnd 7.58fF
C2249 XNOR2X1_11/a_2_6# Gnd 2.31fF
C2250 XNOR2X1_11/a_12_41# Gnd 3.38fF
C2251 XNOR2X1_11/A Gnd 6.68fF
C2252 NAND2X1_13/Y Gnd 11.88fF
C2253 XNOR2X1_24/Y Gnd 9.91fF
C2254 XOR2X1_27/a_2_6# Gnd 3.50fF
C2255 XOR2X1_27/a_13_43# Gnd 3.05fF
C2256 NOR2X1_8/Y Gnd 4.55fF
C2257 INVX2_39/A Gnd 24.04fF
C2258 XNOR2X1_14/a_2_6# Gnd 2.31fF
C2259 XNOR2X1_14/a_12_41# Gnd 3.38fF
C2260 XOR2X1_40/A Gnd 9.01fF
C2261 XOR2X1_29/Y Gnd 5.19fF
C2262 XOR2X1_29/a_2_6# Gnd 3.50fF
C2263 XOR2X1_29/a_13_43# Gnd 3.05fF
C2264 XOR2X1_29/A Gnd 4.27fF
C2265 NOR2X1_9/Y Gnd 5.39fF
C2266 NAND2X1_7/A Gnd 15.82fF
C2267 NOR2X1_9/B Gnd 6.79fF
C2268 XOR2X1_31/a_2_6# Gnd 3.50fF
C2269 XOR2X1_31/a_13_43# Gnd 3.05fF
C2270 NOR2X1_9/A Gnd 9.34fF
C2271 XOR2X1_43/Y Gnd 6.87fF
C2272 XOR2X1_43/B Gnd 11.07fF
C2273 XNOR2X1_16/a_2_6# Gnd 2.31fF
C2274 XNOR2X1_16/a_12_41# Gnd 3.38fF
C2275 INVX2_29/A Gnd 16.51fF
C2276 XOR2X1_81/A Gnd 15.71fF
C2277 XOR2X1_32/Y Gnd 11.65fF
C2278 XOR2X1_32/a_2_6# Gnd 3.50fF
C2279 XOR2X1_32/a_13_43# Gnd 3.05fF
C2280 in_reset Gnd 13.21fF
C2281 XOR2X1_33/B Gnd 13.53fF
C2282 out_MuxData[1] Gnd 18.24fF
C2283 OAI21X1_33/B Gnd 13.45fF
C2284 AOI21X1_4/Y Gnd 7.99fF
C2285 out_state[0] Gnd 17.88fF
C2286 INVX2_31/Y Gnd 10.26fF
C2287 INVX2_34/Y Gnd 10.72fF
C2288 INVX2_32/Y Gnd 6.76fF
C2289 AOI21X1_3/Y Gnd 6.27fF
C2290 DFFPOSX1_16/a_66_6# Gnd 2.23fF
C2291 DFFPOSX1_16/a_2_6# Gnd 3.02fF
C2292 INVX2_36/A Gnd 4.78fF
C2293 AOI22X1_29/C Gnd 3.15fF
C2294 DFFPOSX1_17/a_66_6# Gnd 2.23fF
C2295 DFFPOSX1_17/a_2_6# Gnd 3.02fF
C2296 INVX2_36/Y Gnd 9.35fF
C2297 NAND2X1_10/Y Gnd 5.88fF
C2298 INVX2_44/A Gnd 19.33fF
C2299 DFFPOSX1_18/a_66_6# Gnd 2.23fF
C2300 out_temp_addNum[2] Gnd 22.42fF
C2301 DFFPOSX1_18/a_2_6# Gnd 3.02fF
C2302 OAI21X1_29/Y Gnd 7.50fF
C2303 OR2X2_0/Y Gnd 51.41fF
C2304 DFFPOSX1_23/a_66_6# Gnd 2.23fF
C2305 DFFPOSX1_23/a_2_6# Gnd 3.02fF
C2306 OAI21X1_31/Y Gnd 10.98fF
C2307 XOR2X1_33/a_2_6# Gnd 3.50fF
C2308 XOR2X1_33/a_13_43# Gnd 3.05fF
C2309 AND2X2_15/a_2_6# Gnd 2.37fF
C2310 OAI21X1_32/C Gnd 8.53fF
C2311 XOR2X1_33/A Gnd 7.34fF
C2312 XOR2X1_35/a_2_6# Gnd 3.50fF
C2313 XOR2X1_35/a_13_43# Gnd 3.05fF
C2314 XNOR2X1_17/a_2_6# Gnd 2.31fF
C2315 XNOR2X1_17/a_12_41# Gnd 3.38fF
C2316 XOR2X1_39/Y Gnd 11.52fF
C2317 XOR2X1_39/a_2_6# Gnd 3.50fF
C2318 XOR2X1_39/a_13_43# Gnd 3.05fF
C2319 XOR2X1_40/Y Gnd 9.97fF
C2320 XOR2X1_40/a_2_6# Gnd 3.50fF
C2321 XOR2X1_40/a_13_43# Gnd 3.05fF
C2322 AND2X2_16/Y Gnd 4.04fF
C2323 AND2X2_16/a_2_6# Gnd 2.37fF
C2324 AOI22X1_35/A Gnd 7.43fF
C2325 XNOR2X1_19/a_2_6# Gnd 2.31fF
C2326 XNOR2X1_19/a_12_41# Gnd 3.38fF
C2327 INVX2_86/A Gnd 23.64fF
C2328 XOR2X1_41/a_2_6# Gnd 3.50fF
C2329 XOR2X1_41/a_13_43# Gnd 3.05fF
C2330 XOR2X1_42/a_2_6# Gnd 3.50fF
C2331 XOR2X1_42/a_13_43# Gnd 3.05fF
C2332 XOR2X1_41/A Gnd 4.21fF
C2333 XOR2X1_43/a_2_6# Gnd 3.50fF
C2334 XOR2X1_43/a_13_43# Gnd 3.05fF
C2335 AND2X2_18/A Gnd 8.78fF
C2336 XNOR2X1_21/a_2_6# Gnd 2.31fF
C2337 XNOR2X1_21/a_12_41# Gnd 3.38fF
C2338 XOR2X1_42/A Gnd 5.49fF
C2339 XNOR2X1_22/a_2_6# Gnd 2.31fF
C2340 XNOR2X1_22/a_12_41# Gnd 3.38fF
C2341 XNOR2X1_23/a_2_6# Gnd 2.31fF
C2342 XNOR2X1_23/a_12_41# Gnd 3.38fF
C2343 XOR2X1_50/B Gnd 6.78fF
C2344 NOR2X1_12/B Gnd 11.68fF
C2345 BUFX2_11/Y Gnd 98.79fF
C2346 INVX2_37/Y Gnd 7.13fF
C2347 NOR2X1_14/Y Gnd 14.31fF
C2348 INVX2_50/Y Gnd 42.85fF
C2349 XNOR2X1_27/Y Gnd 6.10fF
C2350 out_MuxData[3] Gnd 35.51fF
C2351 AOI21X1_4/A Gnd 7.84fF
C2352 INVX2_70/Y Gnd 8.08fF
C2353 NAND3X1_12/Y Gnd 9.40fF
C2354 OAI21X1_27/Y Gnd 4.92fF
C2355 NOR2X1_10/B Gnd 11.41fF
C2356 INVX2_35/A Gnd 10.25fF
C2357 NAND2X1_11/Y Gnd 3.88fF
C2358 AOI21X1_5/Y Gnd 8.67fF
C2359 DFFPOSX1_19/a_66_6# Gnd 2.23fF
C2360 DFFPOSX1_19/a_2_6# Gnd 3.02fF
C2361 INVX2_40/A Gnd 13.13fF
C2362 DFFPOSX1_20/a_66_6# Gnd 2.23fF
C2363 DFFPOSX1_20/a_2_6# Gnd 3.02fF
C2364 INVX2_42/Y Gnd 3.63fF
C2365 OAI21X1_38/C Gnd 5.39fF
C2366 DFFPOSX1_21/a_66_6# Gnd 2.23fF
C2367 out_temp_addNum[1] Gnd 27.86fF
C2368 DFFPOSX1_21/a_2_6# Gnd 3.02fF
C2369 OAI21X1_38/Y Gnd 2.71fF
C2370 in_clkb Gnd 68.58fF
C2371 DFFPOSX1_22/a_66_6# Gnd 2.23fF
C2372 DFFPOSX1_22/a_2_6# Gnd 3.02fF
C2373 OAI21X1_30/Y Gnd 8.89fF
C2374 INVX2_38/Y Gnd 7.36fF
C2375 XOR2X1_34/Y Gnd 7.21fF
C2376 XOR2X1_34/a_2_6# Gnd 3.50fF
C2377 XOR2X1_34/a_13_43# Gnd 3.05fF
C2378 XOR2X1_34/A Gnd 12.24fF
C2379 XOR2X1_36/a_2_6# Gnd 3.50fF
C2380 XOR2X1_36/a_13_43# Gnd 3.05fF
C2381 XOR2X1_36/B Gnd 10.56fF
C2382 XOR2X1_37/B Gnd 10.94fF
C2383 XOR2X1_37/a_2_6# Gnd 3.50fF
C2384 XOR2X1_37/a_13_43# Gnd 3.05fF
C2385 NOR2X1_15/B Gnd 5.81fF
C2386 AND2X2_20/Y Gnd 8.56fF
C2387 XNOR2X1_18/a_2_6# Gnd 2.31fF
C2388 XNOR2X1_18/a_12_41# Gnd 3.38fF
C2389 XOR2X1_38/Y Gnd 8.73fF
C2390 XOR2X1_69/B Gnd 48.65fF
C2391 XOR2X1_38/a_2_6# Gnd 3.50fF
C2392 XOR2X1_38/a_13_43# Gnd 3.05fF
C2393 NAND3X1_16/A Gnd 4.93fF
C2394 INVX2_59/Y Gnd 26.91fF
C2395 XNOR2X1_20/a_2_6# Gnd 2.31fF
C2396 XNOR2X1_20/a_12_41# Gnd 3.38fF
C2397 AND2X2_17/Y Gnd 13.51fF
C2398 AND2X2_17/a_2_6# Gnd 2.37fF
C2399 AND2X2_17/B Gnd 3.05fF
C2400 XOR2X1_47/Y Gnd 19.31fF
C2401 XOR2X1_44/Y Gnd 5.27fF
C2402 XOR2X1_44/a_2_6# Gnd 3.50fF
C2403 XOR2X1_44/a_13_43# Gnd 3.05fF
C2404 AND2X2_18/B Gnd 12.92fF
C2405 XNOR2X1_27/A Gnd 6.39fF
C2406 NAND3X1_15/B Gnd 4.47fF
C2407 NAND3X1_15/Y Gnd 9.10fF
C2408 AOI22X1_36/Y Gnd 17.20fF
C2409 BUFX2_3/Y Gnd 20.74fF
C2410 AOI22X1_38/A Gnd 4.76fF
C2411 OAI21X1_39/C Gnd 6.52fF
C2412 INVX2_48/Y Gnd 3.59fF
C2413 XOR2X1_48/B Gnd 11.48fF
C2414 DFFPOSX1_24/a_66_6# Gnd 2.23fF
C2415 DFFPOSX1_24/a_2_6# Gnd 3.02fF
C2416 DFFPOSX1_25/a_66_6# Gnd 2.23fF
C2417 INVX2_52/A Gnd 20.15fF
C2418 DFFPOSX1_25/a_2_6# Gnd 3.02fF
C2419 OAI21X1_35/B Gnd 3.31fF
C2420 INVX2_53/A Gnd 6.62fF
C2421 DFFPOSX1_28/a_66_6# Gnd 2.23fF
C2422 DFFPOSX1_28/a_2_6# Gnd 3.02fF
C2423 INVX2_57/Y Gnd 15.83fF
C2424 INVX2_42/A Gnd 3.03fF
C2425 INVX2_44/Y Gnd 3.59fF
C2426 INVX2_46/A Gnd 24.10fF
C2427 INVX2_47/Y Gnd 5.18fF
C2428 BUFX2_4/Y Gnd 44.86fF
C2429 DFFPOSX1_32/a_66_6# Gnd 2.23fF
C2430 INVX2_48/A Gnd 5.36fF
C2431 DFFPOSX1_32/a_2_6# Gnd 3.02fF
C2432 OAI22X1_1/Y Gnd 4.96fF
C2433 XNOR2X1_24/a_2_6# Gnd 2.31fF
C2434 XNOR2X1_24/a_12_41# Gnd 3.38fF
C2435 NOR2X1_14/A Gnd 11.43fF
C2436 XOR2X1_46/Y Gnd 7.00fF
C2437 XOR2X1_46/a_2_6# Gnd 3.50fF
C2438 XOR2X1_46/a_13_43# Gnd 3.05fF
C2439 OAI21X1_40/A Gnd 12.78fF
C2440 AND2X2_38/Y Gnd 13.51fF
C2441 NOR2X1_15/A Gnd 9.35fF
C2442 AOI22X1_44/Y Gnd 5.31fF
C2443 XNOR2X1_26/a_2_6# Gnd 2.31fF
C2444 XNOR2X1_26/a_12_41# Gnd 3.38fF
C2445 AND2X2_18/a_2_6# Gnd 2.37fF
C2446 XNOR2X1_27/a_2_6# Gnd 2.31fF
C2447 XNOR2X1_27/a_12_41# Gnd 3.38fF
C2448 NOR2X1_17/B Gnd 13.02fF
C2449 XOR2X1_50/Y Gnd 9.81fF
C2450 XOR2X1_50/a_2_6# Gnd 3.50fF
C2451 XOR2X1_50/a_13_43# Gnd 3.05fF
C2452 NOR2X1_13/Y Gnd 2.73fF
C2453 INVX2_62/Y Gnd 33.50fF
C2454 INVX2_87/Y Gnd 37.33fF
C2455 NOR2X1_17/Y Gnd 4.69fF
C2456 DFFPOSX1_26/a_66_6# Gnd 2.23fF
C2457 DFFPOSX1_26/a_2_6# Gnd 3.02fF
C2458 INVX2_40/Y Gnd 14.11fF
C2459 DFFPOSX1_27/a_66_6# Gnd 2.23fF
C2460 INVX2_51/A Gnd 6.47fF
C2461 DFFPOSX1_27/a_2_6# Gnd 3.02fF
C2462 OAI21X1_52/C Gnd 16.54fF
C2463 DFFPOSX1_29/a_66_6# Gnd 2.23fF
C2464 DFFPOSX1_29/a_2_6# Gnd 3.02fF
C2465 OAI21X1_35/Y Gnd 7.11fF
C2466 INVX2_43/Y Gnd 92.52fF
C2467 BUFX2_0/Y Gnd 9.43fF
C2468 BUFX2_0/a_2_6# Gnd 2.75fF
C2469 OAI21X1_44/C Gnd 6.49fF
C2470 con_readData Gnd 40.23fF
C2471 BUFX2_1/Y Gnd 3.83fF
C2472 BUFX2_1/a_2_6# Gnd 2.75fF
C2473 BUFX2_0/A Gnd 9.76fF
C2474 INVX2_46/Y Gnd 14.32fF
C2475 DFFPOSX1_30/a_66_6# Gnd 2.23fF
C2476 out_temp_addNum[0] Gnd 25.91fF
C2477 DFFPOSX1_30/a_2_6# Gnd 3.02fF
C2478 OAI21X1_39/Y Gnd 5.87fF
C2479 DFFPOSX1_31/a_66_6# Gnd 2.23fF
C2480 DFFPOSX1_31/a_2_6# Gnd 3.02fF
C2481 OAI22X1_2/Y Gnd 10.11fF
C2482 INVX2_49/Y Gnd 15.00fF
C2483 INVX2_49/A Gnd 4.67fF
C2484 DFFPOSX1_33/a_66_6# Gnd 2.23fF
C2485 INVX2_65/A Gnd 3.46fF
C2486 DFFPOSX1_33/a_2_6# Gnd 3.02fF
C2487 NOR2X1_14/B Gnd 15.73fF
C2488 XOR2X1_45/a_2_6# Gnd 3.50fF
C2489 XOR2X1_45/a_13_43# Gnd 3.05fF
C2490 XOR2X1_45/Y Gnd 11.33fF
C2491 XNOR2X1_25/a_2_6# Gnd 2.31fF
C2492 XNOR2X1_25/a_12_41# Gnd 3.38fF
C2493 AND2X2_20/B Gnd 5.19fF
C2494 INVX2_92/Y Gnd 17.20fF
C2495 OAI21X1_56/A Gnd 8.46fF
C2496 NOR2X1_16/A Gnd 4.13fF
C2497 INVX2_73/Y Gnd 28.53fF
C2498 XOR2X1_57/Y Gnd 9.49fF
C2499 INVX2_86/Y Gnd 26.34fF
C2500 XOR2X1_47/a_2_6# Gnd 3.50fF
C2501 XOR2X1_47/a_13_43# Gnd 3.05fF
C2502 XOR2X1_52/Y Gnd 9.93fF
C2503 XOR2X1_48/a_2_6# Gnd 3.50fF
C2504 XOR2X1_48/a_13_43# Gnd 3.05fF
C2505 XOR2X1_48/Y Gnd 10.65fF
C2506 XOR2X1_49/Y Gnd 10.02fF
C2507 XOR2X1_49/a_2_6# Gnd 3.50fF
C2508 XOR2X1_49/a_13_43# Gnd 3.05fF
C2509 XOR2X1_49/A Gnd 2.84fF
C2510 OAI21X1_50/B Gnd 11.59fF
C2511 NOR2X1_17/A Gnd 13.40fF
C2512 XNOR2X1_28/a_2_6# Gnd 2.31fF
C2513 XNOR2X1_28/a_12_41# Gnd 3.38fF
C2514 INVX2_56/A Gnd 16.79fF
C2515 NAND2X1_17/B Gnd 7.07fF
C2516 con_writeData Gnd 31.41fF
C2517 OAI21X1_47/C Gnd 4.70fF
C2518 INVX2_65/Y Gnd 8.67fF
C2519 NAND3X1_25/B Gnd 6.31fF
C2520 XOR2X1_55/A Gnd 18.75fF
C2521 AOI22X1_48/Y Gnd 9.20fF
C2522 INVX2_52/Y Gnd 11.23fF
C2523 INVX2_51/Y Gnd 5.86fF
C2524 DFFPOSX1_34/a_66_6# Gnd 2.23fF
C2525 DFFPOSX1_34/a_2_6# Gnd 3.02fF
C2526 INVX2_53/Y Gnd 8.65fF
C2527 OAI21X1_45/C Gnd 5.63fF
C2528 INVX2_54/Y Gnd 9.53fF
C2529 INVX2_58/Y Gnd 9.98fF
C2530 in_DataIn Gnd 16.17fF
C2531 OAI21X1_46/B Gnd 10.36fF
C2532 OR2X2_0/a_2_54# Gnd 2.46fF
C2533 OR2X2_0/B Gnd 6.64fF
C2534 INVX2_59/A Gnd 2.21fF
C2535 out_MemBData[2] Gnd 37.61fF
C2536 INVX2_61/Y Gnd 70.06fF
C2537 DFFPOSX1_37/a_66_6# Gnd 2.23fF
C2538 INVX2_63/A Gnd 7.66fF
C2539 DFFPOSX1_37/a_2_6# Gnd 3.02fF
C2540 OAI22X1_4/Y Gnd 9.85fF
C2541 INVX2_64/Y Gnd 7.71fF
C2542 DFFPOSX1_39/a_66_6# Gnd 2.23fF
C2543 DFFPOSX1_39/a_2_6# Gnd 3.02fF
C2544 INVX2_66/Y Gnd 10.43fF
C2545 INVX2_99/Y Gnd 22.19fF
C2546 INVX2_84/Y Gnd 64.28fF
C2547 DFFPOSX1_40/a_66_6# Gnd 2.23fF
C2548 DFFPOSX1_40/a_2_6# Gnd 3.02fF
C2549 OAI22X1_7/Y Gnd 6.63fF
C2550 AND2X2_20/a_2_6# Gnd 2.37fF
C2551 INVX2_67/Y Gnd 16.36fF
C2552 XNOR2X1_29/a_2_6# Gnd 2.31fF
C2553 XNOR2X1_29/a_12_41# Gnd 3.38fF
C2554 AOI22X1_55/Y Gnd 4.69fF
C2555 XOR2X1_51/a_2_6# Gnd 3.50fF
C2556 XOR2X1_51/a_13_43# Gnd 3.05fF
C2557 XOR2X1_52/a_2_6# Gnd 3.50fF
C2558 XOR2X1_52/a_13_43# Gnd 3.05fF
C2559 XOR2X1_51/Y Gnd 13.09fF
C2560 XNOR2X1_31/a_2_6# Gnd 2.31fF
C2561 XNOR2X1_31/a_12_41# Gnd 3.38fF
C2562 XNOR2X1_32/a_2_6# Gnd 2.31fF
C2563 XNOR2X1_32/a_12_41# Gnd 3.38fF
C2564 XOR2X1_54/A Gnd 19.07fF
C2565 XOR2X1_54/B Gnd 9.52fF
C2566 NAND3X1_22/Y Gnd 3.21fF
C2567 NAND3X1_22/B Gnd 11.42fF
C2568 XOR2X1_53/Y Gnd 4.90fF
C2569 OAI21X1_51/Y Gnd 10.08fF
C2570 INVX2_55/A Gnd 2.98fF
C2571 DFFPOSX1_35/a_66_6# Gnd 2.23fF
C2572 DFFPOSX1_35/a_2_6# Gnd 3.02fF
C2573 INVX2_55/Y Gnd 9.17fF
C2574 INVX2_72/A Gnd 7.03fF
C2575 con_loadData Gnd 25.42fF
C2576 INVX2_57/A Gnd 8.33fF
C2577 OAI21X1_45/Y Gnd 8.16fF
C2578 OAI21X1_45/B Gnd 4.32fF
C2579 AND2X2_19/a_2_6# Gnd 2.37fF
C2580 OR2X2_0/A Gnd 17.82fF
C2581 DFFPOSX1_36/a_66_6# Gnd 2.23fF
C2582 DFFPOSX1_36/a_2_6# Gnd 3.02fF
C2583 OAI21X1_47/Y Gnd 9.33fF
C2584 out_MemBData[0] Gnd 24.28fF
C2585 BUFX2_2/a_2_6# Gnd 2.75fF
C2586 BUFX2_3/a_2_6# Gnd 2.75fF
C2587 BUFX2_4/a_2_6# Gnd 2.75fF
C2588 BUFX2_8/A Gnd 20.11fF
C2589 INVX2_60/Y Gnd 7.41fF
C2590 DFFPOSX1_38/a_66_6# Gnd 2.23fF
C2591 DFFPOSX1_38/a_2_6# Gnd 3.02fF
C2592 INVX2_66/A Gnd 5.75fF
C2593 OAI22X1_6/Y Gnd 6.14fF
C2594 INVX2_63/Y Gnd 20.32fF
C2595 DFFPOSX1_41/a_66_6# Gnd 2.23fF
C2596 DFFPOSX1_41/a_2_6# Gnd 3.02fF
C2597 OAI22X1_8/Y Gnd 9.49fF
C2598 INVX2_67/A Gnd 4.82fF
C2599 AND2X2_23/Y Gnd 9.45fF
C2600 XNOR2X1_30/a_2_6# Gnd 2.31fF
C2601 XNOR2X1_30/a_12_41# Gnd 3.38fF
C2602 OAI21X1_49/Y Gnd 8.41fF
C2603 AND2X2_21/a_2_6# Gnd 2.37fF
C2604 AND2X2_21/A Gnd 9.06fF
C2605 INVX2_94/Y Gnd 24.44fF
C2606 XOR2X1_53/a_2_6# Gnd 3.50fF
C2607 XOR2X1_53/a_13_43# Gnd 3.05fF
C2608 XOR2X1_54/Y Gnd 6.62fF
C2609 XOR2X1_54/a_2_6# Gnd 3.50fF
C2610 XOR2X1_54/a_13_43# Gnd 3.05fF
C2611 AND2X2_22/a_2_6# Gnd 2.37fF
C2612 AOI22X1_48/D Gnd 9.20fF
C2613 AND2X2_22/Y Gnd 3.62fF
C2614 XNOR2X1_33/a_2_6# Gnd 2.31fF
C2615 XNOR2X1_33/a_12_41# Gnd 3.38fF
C2616 AND2X2_24/Y Gnd 6.08fF
C2617 XNOR2X1_34/a_2_6# Gnd 2.31fF
C2618 XNOR2X1_34/a_12_41# Gnd 3.38fF
C2619 OAI21X1_58/Y Gnd 12.43fF
C2620 INVX2_69/A Gnd 5.97fF
C2621 out_MemBData[15] Gnd 35.33fF
C2622 NAND3X1_25/Y Gnd 8.58fF
C2623 XOR2X1_56/Y Gnd 17.81fF
C2624 OAI21X1_59/C Gnd 3.61fF
C2625 DFFPOSX1_43/a_66_6# Gnd 2.23fF
C2626 DFFPOSX1_43/a_2_6# Gnd 3.02fF
C2627 INVX2_69/Y Gnd 14.32fF
C2628 DFFPOSX1_44/a_66_6# Gnd 2.23fF
C2629 DFFPOSX1_44/a_2_6# Gnd 3.02fF
C2630 DFFPOSX1_47/a_66_6# Gnd 2.23fF
C2631 DFFPOSX1_47/a_2_6# Gnd 3.02fF
C2632 OAI21X1_54/Y Gnd 7.94fF
C2633 OAI21X1_55/Y Gnd 3.75fF
C2634 NOR2X1_20/Y Gnd 2.70fF
C2635 BUFX2_7/a_2_6# Gnd 2.75fF
C2636 INVX2_77/A Gnd 9.11fF
C2637 DFFPOSX1_49/a_66_6# Gnd 2.23fF
C2638 DFFPOSX1_49/a_2_6# Gnd 3.02fF
C2639 INVX2_77/Y Gnd 10.28fF
C2640 AOI22X1_50/B Gnd 8.65fF
C2641 DFFPOSX1_51/a_66_6# Gnd 2.23fF
C2642 DFFPOSX1_51/a_2_6# Gnd 3.02fF
C2643 DFFPOSX1_53/a_66_6# Gnd 2.23fF
C2644 DFFPOSX1_53/a_2_6# Gnd 3.02fF
C2645 OAI22X1_9/Y Gnd 9.92fF
C2646 AND2X2_23/a_2_6# Gnd 2.37fF
C2647 INVX2_75/Y Gnd 9.87fF
C2648 XNOR2X1_45/Y Gnd 4.18fF
C2649 XOR2X1_56/a_2_6# Gnd 3.50fF
C2650 XOR2X1_56/a_13_43# Gnd 3.05fF
C2651 XNOR2X1_35/a_2_6# Gnd 2.31fF
C2652 XNOR2X1_35/a_12_41# Gnd 3.38fF
C2653 INVX2_85/Y Gnd 27.31fF
C2654 XOR2X1_58/a_2_6# Gnd 3.50fF
C2655 XOR2X1_58/a_13_43# Gnd 3.05fF
C2656 OAI21X1_57/C Gnd 7.06fF
C2657 NAND2X1_28/Y Gnd 11.71fF
C2658 XOR2X1_58/B Gnd 18.39fF
C2659 AND2X2_24/a_2_6# Gnd 2.37fF
C2660 XOR2X1_58/A Gnd 16.22fF
C2661 OAI21X1_59/B Gnd 7.15fF
C2662 INVX2_126/A Gnd 19.06fF
C2663 NOR2X1_19/Y Gnd 9.15fF
C2664 INVX2_99/A Gnd 45.34fF
C2665 NOR2X1_27/Y Gnd 3.78fF
C2666 AOI21X1_6/B Gnd 16.08fF
C2667 NOR2X1_28/Y Gnd 4.17fF
C2668 out_win Gnd 11.70fF
C2669 DFFPOSX1_42/a_66_6# Gnd 2.23fF
C2670 DFFPOSX1_42/a_2_6# Gnd 3.02fF
C2671 INVX2_79/Y Gnd 8.70fF
C2672 INVX2_72/Y Gnd 22.29fF
C2673 DFFPOSX1_45/a_66_6# Gnd 2.23fF
C2674 con_count[0] Gnd 5.24fF
C2675 DFFPOSX1_45/a_2_6# Gnd 3.02fF
C2676 INVX2_80/Y Gnd 6.29fF
C2677 BUFX2_5/a_2_6# Gnd 2.75fF
C2678 BUFX2_6/a_2_6# Gnd 2.75fF
C2679 in_clka Gnd 7.29fF
C2680 DFFPOSX1_46/a_66_6# Gnd 2.23fF
C2681 DFFPOSX1_46/a_2_6# Gnd 3.02fF
C2682 OAI21X1_60/Y Gnd 9.54fF
C2683 BUFX2_6/Y Gnd 14.65fF
C2684 OAI21X1_60/C Gnd 2.86fF
C2685 DFFPOSX1_48/a_66_6# Gnd 2.23fF
C2686 DFFPOSX1_48/a_2_6# Gnd 3.02fF
C2687 OAI21X1_61/Y Gnd 3.17fF
C2688 INVX2_73/A Gnd 3.37fF
C2689 INVX2_75/A Gnd 15.40fF
C2690 BUFX2_8/a_2_6# Gnd 2.75fF
C2691 out_MemBData[14] Gnd 36.95fF
C2692 INVX2_76/A Gnd 7.25fF
C2693 DFFPOSX1_50/a_66_6# Gnd 2.23fF
C2694 DFFPOSX1_50/a_2_6# Gnd 3.02fF
C2695 INVX2_76/Y Gnd 5.92fF
C2696 AOI22X1_51/B Gnd 3.08fF
C2697 INVX2_78/A Gnd 9.03fF
C2698 DFFPOSX1_52/a_66_6# Gnd 2.23fF
C2699 DFFPOSX1_52/a_2_6# Gnd 3.02fF
C2700 INVX2_78/Y Gnd 9.03fF
C2701 XOR2X1_60/Y Gnd 11.79fF
C2702 NOR2X1_27/A Gnd 11.76fF
C2703 XOR2X1_55/a_2_6# Gnd 3.50fF
C2704 XOR2X1_55/a_13_43# Gnd 3.05fF
C2705 XOR2X1_63/Y Gnd 7.56fF
C2706 XOR2X1_55/Y Gnd 9.37fF
C2707 XOR2X1_57/a_2_6# Gnd 3.50fF
C2708 XOR2X1_57/a_13_43# Gnd 3.05fF
C2709 NOR2X1_28/B Gnd 6.99fF
C2710 XOR2X1_64/B Gnd 5.25fF
C2711 XNOR2X1_36/a_2_6# Gnd 2.31fF
C2712 XNOR2X1_36/a_12_41# Gnd 3.38fF
C2713 XOR2X1_65/A Gnd 6.74fF
C2714 XNOR2X1_41/Y Gnd 11.56fF
C2715 AOI22X1_58/Y Gnd 7.48fF
C2716 AOI22X1_60/C Gnd 9.38fF
C2717 XOR2X1_62/B Gnd 11.91fF
C2718 DFFPOSX1_54/a_66_6# Gnd 2.23fF
C2719 DFFPOSX1_54/a_2_6# Gnd 3.02fF
C2720 OAI21X1_59/Y Gnd 8.78fF
C2721 AOI22X1_59/C Gnd 8.85fF
C2722 INVX2_80/A Gnd 3.42fF
C2723 INVX2_126/Y Gnd 27.32fF
C2724 NOR2X1_35/Y Gnd 23.84fF
C2725 NOR2X1_21/Y Gnd 20.81fF
C2726 NOR2X1_23/Y Gnd 7.12fF
C2727 OAI21X1_62/Y Gnd 5.44fF
C2728 INVX2_81/A Gnd 4.11fF
C2729 out_MemBData[13] Gnd 41.95fF
C2730 DFFPOSX1_59/a_66_6# Gnd 2.23fF
C2731 DFFPOSX1_59/a_2_6# Gnd 3.02fF
C2732 INVX2_81/Y Gnd 8.65fF
C2733 INVX2_83/A Gnd 3.85fF
C2734 AOI22X1_61/B Gnd 9.22fF
C2735 INVX2_83/Y Gnd 5.21fF
C2736 XOR2X1_60/a_2_6# Gnd 3.50fF
C2737 XOR2X1_60/a_13_43# Gnd 3.05fF
C2738 XNOR2X1_37/a_2_6# Gnd 2.31fF
C2739 XNOR2X1_37/a_12_41# Gnd 3.38fF
C2740 XOR2X1_61/a_2_6# Gnd 3.50fF
C2741 XOR2X1_61/a_13_43# Gnd 3.05fF
C2742 XOR2X1_61/Y Gnd 8.90fF
C2743 XNOR2X1_38/a_2_6# Gnd 2.31fF
C2744 XNOR2X1_38/a_12_41# Gnd 3.38fF
C2745 NOR2X1_28/A Gnd 12.85fF
C2746 XOR2X1_64/Y Gnd 7.88fF
C2747 XOR2X1_64/a_2_6# Gnd 3.50fF
C2748 XOR2X1_64/a_13_43# Gnd 3.05fF
C2749 XOR2X1_65/Y Gnd 9.56fF
C2750 XOR2X1_65/a_2_6# Gnd 3.50fF
C2751 XOR2X1_65/a_13_43# Gnd 3.05fF
C2752 NOR2X1_34/Y Gnd 20.32fF
C2753 AOI22X1_62/B Gnd 16.75fF
C2754 DFFPOSX1_55/a_66_6# Gnd 2.23fF
C2755 con_count[7] Gnd 19.19fF
C2756 DFFPOSX1_55/a_2_6# Gnd 3.02fF
C2757 DFFPOSX1_56/a_66_6# Gnd 2.23fF
C2758 DFFPOSX1_56/a_2_6# Gnd 3.02fF
C2759 XOR2X1_59/a_2_6# Gnd 3.50fF
C2760 XOR2X1_59/a_13_43# Gnd 3.05fF
C2761 HAX1_7/YC Gnd 10.44fF
C2762 AND2X2_25/Y Gnd 9.79fF
C2763 AND2X2_25/a_2_6# Gnd 2.37fF
C2764 XOR2X1_59/Y Gnd 2.96fF
C2765 DFFPOSX1_57/a_66_6# Gnd 2.23fF
C2766 DFFPOSX1_57/a_2_6# Gnd 3.02fF
C2767 AND2X2_26/Y Gnd 8.25fF
C2768 AND2X2_26/a_2_6# Gnd 2.37fF
C2769 BUFX2_9/a_2_6# Gnd 2.75fF
C2770 INVX2_91/Y Gnd 15.03fF
C2771 INVX2_90/Y Gnd 13.55fF
C2772 BUFX2_10/a_2_6# Gnd 2.75fF
C2773 DFFPOSX1_58/a_66_6# Gnd 2.23fF
C2774 DFFPOSX1_58/a_2_6# Gnd 3.02fF
C2775 OAI21X1_67/Y Gnd 7.90fF
C2776 OAI21X1_67/C Gnd 5.01fF
C2777 NOR2X1_25/Y Gnd 3.58fF
C2778 INVX2_96/A Gnd 2.43fF
C2779 DFFPOSX1_60/a_66_6# Gnd 2.23fF
C2780 DFFPOSX1_60/a_2_6# Gnd 3.02fF
C2781 INVX2_96/Y Gnd 5.81fF
C2782 INVX2_82/A Gnd 6.02fF
C2783 DFFPOSX1_61/a_66_6# Gnd 2.23fF
C2784 DFFPOSX1_61/a_2_6# Gnd 3.02fF
C2785 INVX2_82/Y Gnd 9.29fF
C2786 DFFPOSX1_62/a_66_6# Gnd 2.23fF
C2787 DFFPOSX1_62/a_2_6# Gnd 3.02fF
C2788 BUFX2_10/Y Gnd 83.06fF
C2789 DFFPOSX1_63/a_66_6# Gnd 2.23fF
C2790 DFFPOSX1_63/a_2_6# Gnd 3.02fF
C2791 INVX2_98/Y Gnd 3.69fF
C2792 XOR2X1_62/Y Gnd 8.31fF
C2793 XOR2X1_62/a_2_6# Gnd 3.50fF
C2794 XOR2X1_62/a_13_43# Gnd 3.05fF
C2795 XOR2X1_63/a_2_6# Gnd 3.50fF
C2796 XOR2X1_63/a_13_43# Gnd 3.05fF
C2797 NAND3X1_27/Y Gnd 4.67fF
C2798 OAI21X1_68/A Gnd 9.33fF
C2799 OAI21X1_68/B Gnd 15.36fF
C2800 XNOR2X1_39/a_2_6# Gnd 2.31fF
C2801 XNOR2X1_39/a_12_41# Gnd 3.38fF
C2802 AND2X2_28/B Gnd 3.68fF
C2803 XNOR2X1_40/a_2_6# Gnd 2.31fF
C2804 XNOR2X1_40/a_12_41# Gnd 3.38fF
C2805 XOR2X1_66/Y Gnd 8.10fF
C2806 XOR2X1_66/a_2_6# Gnd 3.50fF
C2807 XOR2X1_66/a_13_43# Gnd 3.05fF
C2808 XOR2X1_65/B Gnd 8.79fF
C2809 NOR2X1_29/A Gnd 9.85fF
C2810 XNOR2X1_41/a_2_6# Gnd 2.31fF
C2811 XNOR2X1_41/a_12_41# Gnd 3.38fF
C2812 NOR2X1_29/B Gnd 9.23fF
C2813 XOR2X1_74/Y Gnd 16.39fF
C2814 XNOR2X1_42/a_2_6# Gnd 2.31fF
C2815 XNOR2X1_42/a_12_41# Gnd 3.38fF
C2816 INVX2_94/A Gnd 6.59fF
C2817 INVX2_95/Y Gnd 12.33fF
C2818 INVX2_88/A Gnd 5.22fF
C2819 AOI22X1_67/C Gnd 11.40fF
C2820 OR2X1_2/Y Gnd 7.75fF
C2821 OR2X1_2/a_2_54# Gnd 2.68fF
C2822 HAX1_7/YS Gnd 11.70fF
C2823 HAX1_7/a_41_74# Gnd 2.55fF
C2824 HAX1_7/a_2_74# Gnd 2.94fF
C2825 HAX1_7/B Gnd 7.03fF
C2826 AOI22X1_68/C Gnd 9.03fF
C2827 INVX2_89/Y Gnd 7.63fF
C2828 con_count[1] Gnd 39.26fF
C2829 BUFX2_11/a_2_6# Gnd 2.75fF
C2830 INVX2_92/A Gnd 14.28fF
C2831 INVX2_93/A Gnd 16.05fF
C2832 NOR2X1_32/Y Gnd 6.38fF
C2833 DFFPOSX1_69/a_66_6# Gnd 2.23fF
C2834 DFFPOSX1_69/a_2_6# Gnd 3.02fF
C2835 INVX2_97/Y Gnd 8.75fF
C2836 AND2X2_36/A Gnd 15.86fF
C2837 XNOR2X1_43/a_2_6# Gnd 2.31fF
C2838 XNOR2X1_43/a_12_41# Gnd 3.38fF
C2839 XOR2X1_67/a_2_6# Gnd 3.50fF
C2840 XOR2X1_67/a_13_43# Gnd 3.05fF
C2841 AOI21X1_7/B Gnd 16.60fF
C2842 XOR2X1_67/Y Gnd 9.75fF
C2843 XOR2X1_67/B Gnd 9.21fF
C2844 XNOR2X1_44/a_2_6# Gnd 2.31fF
C2845 XNOR2X1_44/a_12_41# Gnd 3.38fF
C2846 XNOR2X1_45/a_2_6# Gnd 2.31fF
C2847 XNOR2X1_45/a_12_41# Gnd 3.38fF
C2848 AND2X2_28/Y Gnd 2.54fF
C2849 AND2X2_28/a_2_6# Gnd 2.37fF
C2850 XNOR2X1_45/A Gnd 5.58fF
C2851 NAND3X1_27/B Gnd 11.47fF
C2852 XOR2X1_72/a_2_6# Gnd 3.50fF
C2853 XOR2X1_72/a_13_43# Gnd 3.05fF
C2854 XOR2X1_72/B Gnd 12.24fF
C2855 XOR2X1_74/B Gnd 13.41fF
C2856 INVX2_95/A Gnd 8.71fF
C2857 OAI22X1_13/Y Gnd 5.79fF
C2858 XOR2X1_69/A Gnd 7.60fF
C2859 DFFPOSX1_64/a_66_6# Gnd 2.23fF
C2860 DFFPOSX1_64/a_2_6# Gnd 3.02fF
C2861 AND2X2_27/Y Gnd 10.12fF
C2862 AND2X2_27/a_2_6# Gnd 2.37fF
C2863 DFFPOSX1_65/a_66_6# Gnd 2.23fF
C2864 DFFPOSX1_65/a_2_6# Gnd 3.02fF
C2865 AND2X2_29/Y Gnd 5.68fF
C2866 DFFPOSX1_66/a_66_6# Gnd 2.23fF
C2867 DFFPOSX1_66/a_2_6# Gnd 3.02fF
C2868 OAI21X1_65/C Gnd 6.80fF
C2869 DFFPOSX1_67/a_66_6# Gnd 2.23fF
C2870 DFFPOSX1_67/a_2_6# Gnd 3.02fF
C2871 OAI21X1_65/Y Gnd 9.85fF
C2872 out_MemBData[4] Gnd 20.96fF
C2873 DFFPOSX1_68/a_66_6# Gnd 2.23fF
C2874 DFFPOSX1_68/a_2_6# Gnd 3.02fF
C2875 INVX2_97/A Gnd 4.77fF
C2876 AOI22X1_69/B Gnd 11.29fF
C2877 INVX2_98/A Gnd 7.82fF
C2878 AOI22X1_80/B Gnd 6.10fF
C2879 DFFPOSX1_70/a_66_6# Gnd 2.23fF
C2880 DFFPOSX1_70/a_2_6# Gnd 3.02fF
C2881 INVX2_109/Y Gnd 9.45fF
C2882 DFFPOSX1_71/a_66_6# Gnd 2.23fF
C2883 DFFPOSX1_71/a_2_6# Gnd 3.02fF
C2884 OAI22X1_10/Y Gnd 8.81fF
C2885 XOR2X1_68/a_2_6# Gnd 3.50fF
C2886 XOR2X1_68/a_13_43# Gnd 3.05fF
C2887 XOR2X1_68/B Gnd 11.62fF
C2888 XOR2X1_69/a_2_6# Gnd 3.50fF
C2889 XOR2X1_69/a_13_43# Gnd 3.05fF
C2890 XOR2X1_70/a_2_6# Gnd 3.50fF
C2891 XOR2X1_70/a_13_43# Gnd 3.05fF
C2892 NOR2X1_42/A Gnd 16.32fF
C2893 XOR2X1_70/B Gnd 5.67fF
C2894 XOR2X1_87/B Gnd 9.71fF
C2895 XOR2X1_70/Y Gnd 11.95fF
C2896 XNOR2X1_46/a_2_6# Gnd 2.31fF
C2897 XNOR2X1_46/a_12_41# Gnd 3.38fF
C2898 XOR2X1_71/a_2_6# Gnd 3.50fF
C2899 XOR2X1_71/a_13_43# Gnd 3.05fF
C2900 OAI21X1_89/A Gnd 13.21fF
C2901 XOR2X1_71/Y Gnd 8.34fF
C2902 XOR2X1_73/a_2_6# Gnd 3.50fF
C2903 XOR2X1_73/a_13_43# Gnd 3.05fF
C2904 XOR2X1_74/a_2_6# Gnd 3.50fF
C2905 XOR2X1_74/a_13_43# Gnd 3.05fF
C2906 con_count[6] Gnd 22.94fF
C2907 NOR2X1_40/Y Gnd 6.55fF
C2908 INVX2_106/A Gnd 11.21fF
C2909 INVX2_107/A Gnd 6.68fF
C2910 AOI22X1_99/Y Gnd 4.47fF
C2911 XOR2X1_90/A Gnd 16.28fF
C2912 DFFPOSX1_72/a_66_6# Gnd 2.23fF
C2913 DFFPOSX1_72/a_2_6# Gnd 3.02fF
C2914 INVX2_102/Y Gnd 8.03fF
C2915 NOR2X1_33/Y Gnd 4.46fF
C2916 AND2X2_29/a_2_6# Gnd 2.37fF
C2917 HAX1_8/YS Gnd 4.95fF
C2918 HAX1_10/B Gnd 11.10fF
C2919 HAX1_8/a_41_74# Gnd 2.55fF
C2920 HAX1_8/a_2_74# Gnd 2.94fF
C2921 AND2X2_30/a_2_6# Gnd 2.37fF
C2922 con_count[2] Gnd 24.64fF
C2923 con_count[3] Gnd 34.36fF
C2924 DFFPOSX1_74/a_66_6# Gnd 2.23fF
C2925 DFFPOSX1_74/a_2_6# Gnd 3.02fF
C2926 OAI21X1_69/Y Gnd 6.29fF
C2927 out_MemBData[9] Gnd 13.89fF
C2928 DFFPOSX1_75/a_66_6# Gnd 2.23fF
C2929 DFFPOSX1_75/a_2_6# Gnd 3.02fF
C2930 INVX2_107/Y Gnd 8.04fF
C2931 INVX2_105/Y Gnd 13.20fF
C2932 DFFPOSX1_76/a_66_6# Gnd 2.23fF
C2933 INVX2_109/A Gnd 5.26fF
C2934 DFFPOSX1_76/a_2_6# Gnd 3.02fF
C2935 OAI22X1_12/Y Gnd 8.60fF
C2936 DFFPOSX1_79/a_66_6# Gnd 2.23fF
C2937 DFFPOSX1_79/a_2_6# Gnd 3.02fF
C2938 OAI22X1_14/Y Gnd 7.42fF
C2939 AOI21X1_7/A Gnd 15.20fF
C2940 XNOR2X1_47/a_2_6# Gnd 2.31fF
C2941 XNOR2X1_47/a_12_41# Gnd 3.38fF
C2942 XOR2X1_75/Y Gnd 14.00fF
C2943 XOR2X1_75/a_2_6# Gnd 3.50fF
C2944 XOR2X1_75/a_13_43# Gnd 3.05fF
C2945 XOR2X1_76/Y Gnd 8.08fF
C2946 XOR2X1_76/a_2_6# Gnd 3.50fF
C2947 XOR2X1_76/a_13_43# Gnd 3.05fF
C2948 AOI22X1_96/Y Gnd 9.12fF
C2949 XNOR2X1_49/a_2_6# Gnd 2.31fF
C2950 XNOR2X1_49/a_12_41# Gnd 3.38fF
C2951 XOR2X1_80/a_2_6# Gnd 3.50fF
C2952 XOR2X1_80/a_13_43# Gnd 3.05fF
C2953 NOR2X1_45/A Gnd 10.45fF
C2954 XOR2X1_84/B Gnd 7.79fF
C2955 INVX2_120/A Gnd 15.42fF
C2956 OAI21X1_71/Y Gnd 10.73fF
C2957 out_MemBData[5] Gnd 23.37fF
C2958 OAI21X1_73/Y Gnd 3.82fF
C2959 INVX2_102/A Gnd 6.87fF
C2960 DFFPOSX1_73/a_66_6# Gnd 2.23fF
C2961 AOI22X1_79/C Gnd 2.31fF
C2962 DFFPOSX1_73/a_2_6# Gnd 3.02fF
C2963 HAX1_9/a_41_74# Gnd 2.55fF
C2964 HAX1_9/a_2_74# Gnd 2.94fF
C2965 HAX1_9/B Gnd 7.25fF
C2966 AND2X2_31/Y Gnd 8.97fF
C2967 AND2X2_31/a_2_6# Gnd 2.37fF
C2968 HAX1_9/YS Gnd 5.17fF
C2969 HAX1_13/B Gnd 12.02fF
C2970 HAX1_10/a_41_74# Gnd 2.55fF
C2971 HAX1_10/a_2_74# Gnd 2.94fF
C2972 NOR2X1_39/A Gnd 7.26fF
C2973 INVX2_103/Y Gnd 12.92fF
C2974 NOR2X1_36/Y Gnd 23.07fF
C2975 INVX2_104/A Gnd 15.73fF
C2976 OAI21X1_71/C Gnd 6.17fF
C2977 out_MemBData[8] Gnd 24.81fF
C2978 NOR2X1_37/Y Gnd 4.96fF
C2979 OAI21X1_73/C Gnd 7.07fF
C2980 NOR2X1_38/Y Gnd 7.40fF
C2981 out_MemBData[10] Gnd 23.14fF
C2982 INVX2_108/Y Gnd 3.31fF
C2983 DFFPOSX1_77/a_66_6# Gnd 2.23fF
C2984 DFFPOSX1_77/a_2_6# Gnd 3.02fF
C2985 OAI22X1_11/Y Gnd 9.14fF
C2986 INVX2_110/A Gnd 4.67fF
C2987 DFFPOSX1_78/a_66_6# Gnd 2.23fF
C2988 DFFPOSX1_78/a_2_6# Gnd 3.02fF
C2989 OAI22X1_16/Y Gnd 7.50fF
C2990 NOR2X1_42/B Gnd 12.67fF
C2991 OAI21X1_78/A Gnd 13.77fF
C2992 XNOR2X1_48/a_2_6# Gnd 2.31fF
C2993 XNOR2X1_48/a_12_41# Gnd 3.38fF
C2994 XOR2X1_77/Y Gnd 11.22fF
C2995 XOR2X1_77/a_2_6# Gnd 3.50fF
C2996 XOR2X1_77/a_13_43# Gnd 3.05fF
C2997 NOR2X1_44/A Gnd 8.23fF
C2998 XOR2X1_78/Y Gnd 7.76fF
C2999 XOR2X1_78/B Gnd 10.59fF
C3000 XOR2X1_78/a_2_6# Gnd 3.50fF
C3001 XOR2X1_78/a_13_43# Gnd 3.05fF
C3002 OAI21X1_91/A Gnd 14.07fF
C3003 XOR2X1_79/Y Gnd 3.07fF
C3004 XOR2X1_79/a_2_6# Gnd 3.50fF
C3005 XOR2X1_79/a_13_43# Gnd 3.05fF
C3006 INVX2_118/A Gnd 16.00fF
C3007 INVX2_130/A Gnd 17.02fF
C3008 INVX2_121/Y Gnd 21.28fF
C3009 NOR2X1_44/B Gnd 14.26fF
C3010 AND2X2_40/A Gnd 13.40fF
C3011 DFFPOSX1_80/a_66_6# Gnd 2.23fF
C3012 AOI22X1_87/C Gnd 8.49fF
C3013 DFFPOSX1_80/a_2_6# Gnd 3.02fF
C3014 HAX1_11/a_41_74# Gnd 2.55fF
C3015 HAX1_11/a_2_74# Gnd 2.94fF
C3016 HAX1_11/B Gnd 9.71fF
C3017 AND2X2_32/Y Gnd 8.71fF
C3018 AND2X2_32/a_2_6# Gnd 2.37fF
C3019 AND2X2_33/a_2_6# Gnd 2.37fF
C3020 DFFPOSX1_81/a_66_6# Gnd 2.23fF
C3021 AOI22X1_88/C Gnd 10.79fF
C3022 DFFPOSX1_81/a_2_6# Gnd 3.02fF
C3023 AND2X2_33/Y Gnd 9.67fF
C3024 INVX2_117/A Gnd 10.34fF
C3025 INVX2_128/A Gnd 7.21fF
C3026 NOR2X1_39/Y Gnd 12.76fF
C3027 DFFPOSX1_83/a_66_6# Gnd 2.23fF
C3028 DFFPOSX1_83/a_2_6# Gnd 3.02fF
C3029 DFFPOSX1_86/a_66_6# Gnd 2.23fF
C3030 DFFPOSX1_86/a_2_6# Gnd 3.02fF
C3031 INVX2_119/Y Gnd 11.57fF
C3032 DFFPOSX1_88/a_66_6# Gnd 2.23fF
C3033 INVX2_121/A Gnd 3.00fF
C3034 DFFPOSX1_88/a_2_6# Gnd 3.02fF
C3035 OAI22X1_15/Y Gnd 7.57fF
C3036 DFFPOSX1_89/a_66_6# Gnd 2.23fF
C3037 DFFPOSX1_89/a_2_6# Gnd 3.02fF
C3038 OAI22X1_18/Y Gnd 2.55fF
C3039 AND2X2_36/B Gnd 12.55fF
C3040 XNOR2X1_50/a_2_6# Gnd 2.31fF
C3041 XNOR2X1_50/a_12_41# Gnd 3.38fF
C3042 OAI21X1_87/A Gnd 22.05fF
C3043 XOR2X1_81/Y Gnd 7.79fF
C3044 XOR2X1_81/a_2_6# Gnd 3.50fF
C3045 XOR2X1_81/a_13_43# Gnd 3.05fF
C3046 XOR2X1_82/B Gnd 5.33fF
C3047 XNOR2X1_51/a_2_6# Gnd 2.31fF
C3048 XNOR2X1_51/a_12_41# Gnd 3.38fF
C3049 OAI21X1_79/C Gnd 11.55fF
C3050 OAI21X1_78/B Gnd 10.87fF
C3051 XOR2X1_87/A Gnd 6.12fF
C3052 XNOR2X1_52/a_2_6# Gnd 2.31fF
C3053 XNOR2X1_52/a_12_41# Gnd 3.38fF
C3054 OAI21X1_89/B Gnd 19.45fF
C3055 XNOR2X1_53/a_2_6# Gnd 2.31fF
C3056 XNOR2X1_53/a_12_41# Gnd 3.38fF
C3057 XNOR2X1_54/a_2_6# Gnd 2.31fF
C3058 XNOR2X1_54/a_12_41# Gnd 3.38fF
C3059 XOR2X1_91/A Gnd 14.45fF
C3060 XNOR2X1_55/a_2_6# Gnd 2.31fF
C3061 XNOR2X1_55/a_12_41# Gnd 3.38fF
C3062 XOR2X1_83/a_2_6# Gnd 3.50fF
C3063 XOR2X1_83/a_13_43# Gnd 3.05fF
C3064 NOR2X1_45/B Gnd 10.43fF
C3065 XOR2X1_83/Y Gnd 10.50fF
C3066 XOR2X1_83/B Gnd 8.15fF
C3067 XOR2X1_84/a_2_6# Gnd 3.50fF
C3068 XOR2X1_84/a_13_43# Gnd 3.05fF
C3069 INVX2_122/A Gnd 9.89fF
C3070 XOR2X1_89/Y Gnd 6.68fF
C3071 INVX2_124/A Gnd 8.01fF
C3072 HAX1_12/a_41_74# Gnd 2.55fF
C3073 HAX1_12/a_2_74# Gnd 2.94fF
C3074 con_count[4] Gnd 19.82fF
C3075 con_count[5] Gnd 21.72fF
C3076 HAX1_12/B Gnd 7.26fF
C3077 HAX1_13/a_41_74# Gnd 2.55fF
C3078 HAX1_13/a_2_74# Gnd 2.94fF
C3079 DFFPOSX1_82/a_66_6# Gnd 2.23fF
C3080 DFFPOSX1_82/a_2_6# Gnd 3.02fF
C3081 INVX2_116/Y Gnd 11.13fF
C3082 INVX2_116/A Gnd 7.25fF
C3083 OAI21X1_81/Y Gnd 7.88fF
C3084 DFFPOSX1_84/a_66_6# Gnd 2.23fF
C3085 DFFPOSX1_84/a_2_6# Gnd 3.02fF
C3086 OAI21X1_75/Y Gnd 8.86fF
C3087 DFFPOSX1_85/a_66_6# Gnd 2.23fF
C3088 DFFPOSX1_85/a_2_6# Gnd 3.02fF
C3089 OAI21X1_83/Y Gnd 3.98fF
C3090 OAI21X1_76/C Gnd 5.33fF
C3091 NOR2X1_41/Y Gnd 5.38fF
C3092 DFFPOSX1_87/a_66_6# Gnd 2.23fF
C3093 out_MemBData[11] Gnd 8.40fF
C3094 DFFPOSX1_87/a_2_6# Gnd 3.02fF
C3095 OAI21X1_76/Y Gnd 14.67fF
C3096 INVX2_133/Y Gnd 12.96fF
C3097 OAI22X1_17/Y Gnd 6.07fF
C3098 INVX2_122/Y Gnd 18.26fF
C3099 INVX2_123/Y Gnd 14.87fF
C3100 INVX2_123/A Gnd 4.47fF
C3101 XOR2X1_85/B Gnd 2.86fF
C3102 XOR2X1_82/Y Gnd 5.44fF
C3103 XOR2X1_82/a_2_6# Gnd 3.50fF
C3104 XOR2X1_82/a_13_43# Gnd 3.05fF
C3105 XOR2X1_82/A Gnd 5.54fF
C3106 OAI21X1_78/C Gnd 6.60fF
C3107 AND2X2_39/B Gnd 4.37fF
C3108 NOR2X1_46/B Gnd 10.46fF
C3109 XOR2X1_88/Y Gnd 6.56fF
C3110 OAI21X1_89/C Gnd 5.39fF
C3111 OAI21X1_90/C Gnd 8.31fF
C3112 AND2X2_41/A Gnd 10.26fF
C3113 XNOR2X1_56/a_2_6# Gnd 2.31fF
C3114 XNOR2X1_56/a_12_41# Gnd 3.38fF
C3115 XOR2X1_89/B Gnd 13.18fF
C3116 AOI22X1_93/C Gnd 3.52fF
C3117 XOR2X1_89/A Gnd 6.42fF
C3118 DFFPOSX1_90/a_66_6# Gnd 2.23fF
C3119 DFFPOSX1_90/a_2_6# Gnd 3.02fF
C3120 INVX2_124/Y Gnd 8.04fF
C3121 AND2X2_34/Y Gnd 7.99fF
C3122 AND2X2_34/a_2_6# Gnd 2.37fF
C3123 INVX2_125/A Gnd 11.63fF
C3124 AND2X2_35/a_2_6# Gnd 2.37fF
C3125 INVX2_127/A Gnd 8.80fF
C3126 DFFPOSX1_93/a_66_6# Gnd 2.23fF
C3127 AOI22X1_94/C Gnd 4.23fF
C3128 DFFPOSX1_93/a_2_6# Gnd 3.02fF
C3129 AND2X2_35/Y Gnd 9.27fF
C3130 NOR2X1_46/Y Gnd 5.42fF
C3131 OAI21X1_84/Y Gnd 2.59fF
C3132 NOR2X1_48/Y Gnd 2.16fF
C3133 DFFPOSX1_96/a_66_6# Gnd 2.23fF
C3134 out_MemBData[7] Gnd 16.54fF
C3135 DFFPOSX1_96/a_2_6# Gnd 3.02fF
C3136 OAI21X1_85/Y Gnd 8.16fF
C3137 INVX2_132/Y Gnd 7.53fF
C3138 DFFPOSX1_97/a_66_6# Gnd 2.23fF
C3139 DFFPOSX1_97/a_2_6# Gnd 3.02fF
C3140 OAI22X1_20/Y Gnd 8.18fF
C3141 DFFPOSX1_98/a_66_6# Gnd 2.23fF
C3142 DFFPOSX1_98/a_2_6# Gnd 3.02fF
C3143 NAND2X1_42/Y Gnd 10.07fF
C3144 XOR2X1_85/a_2_6# Gnd 3.50fF
C3145 XOR2X1_85/a_13_43# Gnd 3.05fF
C3146 XOR2X1_85/A Gnd 7.38fF
C3147 XOR2X1_85/Y Gnd 4.74fF
C3148 NOR2X1_49/B Gnd 15.82fF
C3149 XNOR2X1_58/a_2_6# Gnd 2.31fF
C3150 XNOR2X1_58/a_12_41# Gnd 3.38fF
C3151 AND2X2_37/Y Gnd 6.47fF
C3152 AND2X2_37/a_2_6# Gnd 2.37fF
C3153 AND2X2_39/a_2_6# Gnd 2.37fF
C3154 XOR2X1_88/a_2_6# Gnd 3.50fF
C3155 XOR2X1_88/a_13_43# Gnd 3.05fF
C3156 XOR2X1_88/A Gnd 5.00fF
C3157 AND2X2_40/Y Gnd 6.57fF
C3158 AND2X2_40/a_2_6# Gnd 2.37fF
C3159 AND2X2_41/a_2_6# Gnd 2.37fF
C3160 XOR2X1_89/a_2_6# Gnd 3.50fF
C3161 XOR2X1_89/a_13_43# Gnd 3.05fF
C3162 NAND3X1_34/Y Gnd 5.78fF
C3163 INVX2_135/Y Gnd 14.34fF
C3164 DFFPOSX1_91/a_66_6# Gnd 2.23fF
C3165 DFFPOSX1_91/a_2_6# Gnd 3.02fF
C3166 INVX2_125/Y Gnd 8.19fF
C3167 DFFPOSX1_92/a_66_6# Gnd 2.23fF
C3168 DFFPOSX1_92/a_2_6# Gnd 3.02fF
C3169 DFFPOSX1_94/a_66_6# Gnd 2.23fF
C3170 DFFPOSX1_94/a_2_6# Gnd 3.02fF
C3171 INVX2_127/Y Gnd 8.39fF
C3172 DFFPOSX1_95/a_66_6# Gnd 2.23fF
C3173 DFFPOSX1_95/a_2_6# Gnd 3.02fF
C3174 OAI21X1_80/Y Gnd 9.93fF
C3175 OAI21X1_80/C Gnd 2.09fF
C3176 NOR2X1_47/Y Gnd 5.81fF
C3177 NOR2X1_49/Y Gnd 4.24fF
C3178 INVX2_129/Y Gnd 13.04fF
C3179 INVX2_131/Y Gnd 5.05fF
C3180 DFFPOSX1_99/a_66_6# Gnd 2.23fF
C3181 INVX2_133/A Gnd 10.08fF
C3182 DFFPOSX1_99/a_2_6# Gnd 3.02fF
C3183 OAI22X1_21/Y Gnd 9.33fF
C3184 DFFPOSX1_100/a_66_6# Gnd 2.23fF
C3185 DFFPOSX1_100/a_2_6# Gnd 3.02fF
C3186 OAI22X1_19/Y Gnd 9.20fF
C3187 INVX2_134/A Gnd 5.36fF
C3188 XNOR2X1_57/a_2_6# Gnd 2.31fF
C3189 XNOR2X1_57/a_12_41# Gnd 3.38fF
C3190 OAI21X1_88/Y Gnd 6.26fF
C3191 AND2X2_36/Y Gnd 4.10fF
C3192 AND2X2_36/a_2_6# Gnd 2.37fF
C3193 XOR2X1_86/a_2_6# Gnd 3.50fF
C3194 XOR2X1_86/a_13_43# Gnd 3.05fF
C3195 XNOR2X1_57/Y Gnd 9.64fF
C3196 XOR2X1_86/Y Gnd 4.74fF
C3197 AND2X2_38/a_2_6# Gnd 2.37fF
C3198 AND2X2_38/A Gnd 7.50fF
C3199 XOR2X1_87/Y Gnd 9.06fF
C3200 XOR2X1_87/a_2_6# Gnd 3.50fF
C3201 XOR2X1_87/a_13_43# Gnd 3.05fF
C3202 AND2X2_38/B Gnd 8.19fF
C3203 XOR2X1_90/a_2_6# Gnd 3.50fF
C3204 XOR2X1_90/a_13_43# Gnd 3.05fF
C3205 AOI22X1_99/D Gnd 11.07fF
C3206 XNOR2X1_59/a_2_6# Gnd 2.31fF
C3207 XNOR2X1_59/a_12_41# Gnd 3.38fF
C3208 OAI21X1_90/Y Gnd 9.53fF
C3209 XOR2X1_91/a_2_6# Gnd 3.50fF
C3210 XOR2X1_91/a_13_43# Gnd 3.05fF
C3211 AOI22X1_99/B Gnd 8.55fF
C3212 XNOR2X1_60/a_2_6# Gnd 2.31fF
C3213 XNOR2X1_60/a_12_41# Gnd 3.38fF
C3214 XNOR2X1_60/A Gnd 6.68fF
